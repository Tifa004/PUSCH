module Twiddle960 #(
    parameter   TW_FF = 0   //  Use Output Register
)(
    input           clk,  //  Master Clock
    input   [10:0]   addr,   //  Twiddle Factor Number
    output  [17:0]  tw_re,  //  Twiddle Factor (Real)
    output  [17:0]  tw_im   //  Twiddle Factor (Imag)
);

wire[17:0]  wn_re[0:959];   //  Twiddle Table (Real)
wire[17:0]  wn_im[0:959];   //  Twiddle Table (Imag)
wire[17:0]  mx_re;          //  Multiplexer output (Real)
wire[17:0]  mx_im;          //  Multiplexer output (Imag)
reg [17:0]  ff_re;          //  Register output (Real)
reg [17:0]  ff_im;          //  Register output (Imag)

assign  mx_re = addr<960 ? wn_re[addr] : 0;
assign  mx_im = addr<960 ? wn_im[addr] : 0;

always @(posedge clk) begin
    ff_re <= mx_re;
    ff_im <= mx_im;
end

assign  tw_re = TW_FF ? ff_re : mx_re;
assign  tw_im = TW_FF ? ff_im : mx_im;
assign wn_re[0] = 18'b000000010000000000; assign wn_im[0] = 18'b000000000000000000; 
assign wn_re[1] = 18'b000000001111111111; assign wn_im[1] = 18'b111111111111111001; 
assign wn_re[2] = 18'b000000001111111111; assign wn_im[2] = 18'b111111111111110010; 
assign wn_re[3] = 18'b000000001111111111; assign wn_im[3] = 18'b111111111111101011; 
assign wn_re[4] = 18'b000000001111111111; assign wn_im[4] = 18'b111111111111100101; 
assign wn_re[5] = 18'b000000001111111111; assign wn_im[5] = 18'b111111111111011110; 
assign wn_re[6] = 18'b000000001111111111; assign wn_im[6] = 18'b111111111111010111; 
assign wn_re[7] = 18'b000000001111111110; assign wn_im[7] = 18'b111111111111010001; 
assign wn_re[8] = 18'b000000001111111110; assign wn_im[8] = 18'b111111111111001010; 
assign wn_re[9] = 18'b000000001111111110; assign wn_im[9] = 18'b111111111111000011; 
assign wn_re[10] = 18'b000000001111111101; assign wn_im[10] = 18'b111111111110111101; 
assign wn_re[11] = 18'b000000001111111101; assign wn_im[11] = 18'b111111111110110110; 
assign wn_re[12] = 18'b000000001111111100; assign wn_im[12] = 18'b111111111110101111; 
assign wn_re[13] = 18'b000000001111111100; assign wn_im[13] = 18'b111111111110101000; 
assign wn_re[14] = 18'b000000001111111011; assign wn_im[14] = 18'b111111111110100010; 
assign wn_re[15] = 18'b000000001111111011; assign wn_im[15] = 18'b111111111110011011; 
assign wn_re[16] = 18'b000000001111111010; assign wn_im[16] = 18'b111111111110010100; 
assign wn_re[17] = 18'b000000001111111001; assign wn_im[17] = 18'b111111111110001110; 
assign wn_re[18] = 18'b000000001111111000; assign wn_im[18] = 18'b111111111110000111; 
assign wn_re[19] = 18'b000000001111111000; assign wn_im[19] = 18'b111111111110000000; 
assign wn_re[20] = 18'b000000001111110111; assign wn_im[20] = 18'b111111111101111010; 
assign wn_re[21] = 18'b000000001111110110; assign wn_im[21] = 18'b111111111101110011; 
assign wn_re[22] = 18'b000000001111110101; assign wn_im[22] = 18'b111111111101101101; 
assign wn_re[23] = 18'b000000001111110100; assign wn_im[23] = 18'b111111111101100110; 
assign wn_re[24] = 18'b000000001111110011; assign wn_im[24] = 18'b111111111101011111; 
assign wn_re[25] = 18'b000000001111110010; assign wn_im[25] = 18'b111111111101011001; 
assign wn_re[26] = 18'b000000001111110001; assign wn_im[26] = 18'b111111111101010010; 
assign wn_re[27] = 18'b000000001111110000; assign wn_im[27] = 18'b111111111101001011; 
assign wn_re[28] = 18'b000000001111101110; assign wn_im[28] = 18'b111111111101000101; 
assign wn_re[29] = 18'b000000001111101101; assign wn_im[29] = 18'b111111111100111110; 
assign wn_re[30] = 18'b000000001111101100; assign wn_im[30] = 18'b111111111100111000; 
assign wn_re[31] = 18'b000000001111101010; assign wn_im[31] = 18'b111111111100110001; 
assign wn_re[32] = 18'b000000001111101001; assign wn_im[32] = 18'b111111111100101011; 
assign wn_re[33] = 18'b000000001111101000; assign wn_im[33] = 18'b111111111100100100; 
assign wn_re[34] = 18'b000000001111100110; assign wn_im[34] = 18'b111111111100011110; 
assign wn_re[35] = 18'b000000001111100101; assign wn_im[35] = 18'b111111111100010111; 
assign wn_re[36] = 18'b000000001111100011; assign wn_im[36] = 18'b111111111100010000; 
assign wn_re[37] = 18'b000000001111100010; assign wn_im[37] = 18'b111111111100001010; 
assign wn_re[38] = 18'b000000001111100000; assign wn_im[38] = 18'b111111111100000011; 
assign wn_re[39] = 18'b000000001111011110; assign wn_im[39] = 18'b111111111011111101; 
assign wn_re[40] = 18'b000000001111011101; assign wn_im[40] = 18'b111111111011110110; 
assign wn_re[41] = 18'b000000001111011011; assign wn_im[41] = 18'b111111111011110000; 
assign wn_re[42] = 18'b000000001111011001; assign wn_im[42] = 18'b111111111011101010; 
assign wn_re[43] = 18'b000000001111010111; assign wn_im[43] = 18'b111111111011100011; 
assign wn_re[44] = 18'b000000001111010101; assign wn_im[44] = 18'b111111111011011101; 
assign wn_re[45] = 18'b000000001111010011; assign wn_im[45] = 18'b111111111011010110; 
assign wn_re[46] = 18'b000000001111010001; assign wn_im[46] = 18'b111111111011010000; 
assign wn_re[47] = 18'b000000001111001111; assign wn_im[47] = 18'b111111111011001001; 
assign wn_re[48] = 18'b000000001111001101; assign wn_im[48] = 18'b111111111011000011; 
assign wn_re[49] = 18'b000000001111001011; assign wn_im[49] = 18'b111111111010111101; 
assign wn_re[50] = 18'b000000001111001001; assign wn_im[50] = 18'b111111111010110110; 
assign wn_re[51] = 18'b000000001111000111; assign wn_im[51] = 18'b111111111010110000; 
assign wn_re[52] = 18'b000000001111000101; assign wn_im[52] = 18'b111111111010101010; 
assign wn_re[53] = 18'b000000001111000011; assign wn_im[53] = 18'b111111111010100011; 
assign wn_re[54] = 18'b000000001111000000; assign wn_im[54] = 18'b111111111010011101; 
assign wn_re[55] = 18'b000000001110111110; assign wn_im[55] = 18'b111111111010010111; 
assign wn_re[56] = 18'b000000001110111011; assign wn_im[56] = 18'b111111111010010001; 
assign wn_re[57] = 18'b000000001110111001; assign wn_im[57] = 18'b111111111010001010; 
assign wn_re[58] = 18'b000000001110110111; assign wn_im[58] = 18'b111111111010000100; 
assign wn_re[59] = 18'b000000001110110100; assign wn_im[59] = 18'b111111111001111110; 
assign wn_re[60] = 18'b000000001110110010; assign wn_im[60] = 18'b111111111001111000; 
assign wn_re[61] = 18'b000000001110101111; assign wn_im[61] = 18'b111111111001110001; 
assign wn_re[62] = 18'b000000001110101100; assign wn_im[62] = 18'b111111111001101011; 
assign wn_re[63] = 18'b000000001110101010; assign wn_im[63] = 18'b111111111001100101; 
assign wn_re[64] = 18'b000000001110100111; assign wn_im[64] = 18'b111111111001011111; 
assign wn_re[65] = 18'b000000001110100100; assign wn_im[65] = 18'b111111111001011001; 
assign wn_re[66] = 18'b000000001110100001; assign wn_im[66] = 18'b111111111001010011; 
assign wn_re[67] = 18'b000000001110011111; assign wn_im[67] = 18'b111111111001001101; 
assign wn_re[68] = 18'b000000001110011100; assign wn_im[68] = 18'b111111111001000111; 
assign wn_re[69] = 18'b000000001110011001; assign wn_im[69] = 18'b111111111001000001; 
assign wn_re[70] = 18'b000000001110010110; assign wn_im[70] = 18'b111111111000111011; 
assign wn_re[71] = 18'b000000001110010011; assign wn_im[71] = 18'b111111111000110101; 
assign wn_re[72] = 18'b000000001110010000; assign wn_im[72] = 18'b111111111000101111; 
assign wn_re[73] = 18'b000000001110001101; assign wn_im[73] = 18'b111111111000101001; 
assign wn_re[74] = 18'b000000001110001010; assign wn_im[74] = 18'b111111111000100011; 
assign wn_re[75] = 18'b000000001110000111; assign wn_im[75] = 18'b111111111000011101; 
assign wn_re[76] = 18'b000000001110000011; assign wn_im[76] = 18'b111111111000010111; 
assign wn_re[77] = 18'b000000001110000000; assign wn_im[77] = 18'b111111111000010001; 
assign wn_re[78] = 18'b000000001101111101; assign wn_im[78] = 18'b111111111000001011; 
assign wn_re[79] = 18'b000000001101111010; assign wn_im[79] = 18'b111111111000000101; 
assign wn_re[80] = 18'b000000001101110110; assign wn_im[80] = 18'b111111111000000000; 
assign wn_re[81] = 18'b000000001101110011; assign wn_im[81] = 18'b111111110111111010; 
assign wn_re[82] = 18'b000000001101110000; assign wn_im[82] = 18'b111111110111110100; 
assign wn_re[83] = 18'b000000001101101100; assign wn_im[83] = 18'b111111110111101110; 
assign wn_re[84] = 18'b000000001101101001; assign wn_im[84] = 18'b111111110111101000; 
assign wn_re[85] = 18'b000000001101100101; assign wn_im[85] = 18'b111111110111100011; 
assign wn_re[86] = 18'b000000001101100010; assign wn_im[86] = 18'b111111110111011101; 
assign wn_re[87] = 18'b000000001101011110; assign wn_im[87] = 18'b111111110111010111; 
assign wn_re[88] = 18'b000000001101011010; assign wn_im[88] = 18'b111111110111010010; 
assign wn_re[89] = 18'b000000001101010111; assign wn_im[89] = 18'b111111110111001100; 
assign wn_re[90] = 18'b000000001101010011; assign wn_im[90] = 18'b111111110111000111; 
assign wn_re[91] = 18'b000000001101001111; assign wn_im[91] = 18'b111111110111000001; 
assign wn_re[92] = 18'b000000001101001011; assign wn_im[92] = 18'b111111110110111100; 
assign wn_re[93] = 18'b000000001101001000; assign wn_im[93] = 18'b111111110110110110; 
assign wn_re[94] = 18'b000000001101000100; assign wn_im[94] = 18'b111111110110110001; 
assign wn_re[95] = 18'b000000001101000000; assign wn_im[95] = 18'b111111110110101011; 
assign wn_re[96] = 18'b000000001100111100; assign wn_im[96] = 18'b111111110110100110; 
assign wn_re[97] = 18'b000000001100111000; assign wn_im[97] = 18'b111111110110100000; 
assign wn_re[98] = 18'b000000001100110100; assign wn_im[98] = 18'b111111110110011011; 
assign wn_re[99] = 18'b000000001100110000; assign wn_im[99] = 18'b111111110110010101; 
assign wn_re[100] = 18'b000000001100101100; assign wn_im[100] = 18'b111111110110010000; 
assign wn_re[101] = 18'b000000001100101000; assign wn_im[101] = 18'b111111110110001011; 
assign wn_re[102] = 18'b000000001100100100; assign wn_im[102] = 18'b111111110110000110; 
assign wn_re[103] = 18'b000000001100011111; assign wn_im[103] = 18'b111111110110000000; 
assign wn_re[104] = 18'b000000001100011011; assign wn_im[104] = 18'b111111110101111011; 
assign wn_re[105] = 18'b000000001100010111; assign wn_im[105] = 18'b111111110101110110; 
assign wn_re[106] = 18'b000000001100010011; assign wn_im[106] = 18'b111111110101110001; 
assign wn_re[107] = 18'b000000001100001110; assign wn_im[107] = 18'b111111110101101100; 
assign wn_re[108] = 18'b000000001100001010; assign wn_im[108] = 18'b111111110101100110; 
assign wn_re[109] = 18'b000000001100000110; assign wn_im[109] = 18'b111111110101100001; 
assign wn_re[110] = 18'b000000001100000001; assign wn_im[110] = 18'b111111110101011100; 
assign wn_re[111] = 18'b000000001011111101; assign wn_im[111] = 18'b111111110101010111; 
assign wn_re[112] = 18'b000000001011111000; assign wn_im[112] = 18'b111111110101010010; 
assign wn_re[113] = 18'b000000001011110100; assign wn_im[113] = 18'b111111110101001101; 
assign wn_re[114] = 18'b000000001011101111; assign wn_im[114] = 18'b111111110101001000; 
assign wn_re[115] = 18'b000000001011101011; assign wn_im[115] = 18'b111111110101000100; 
assign wn_re[116] = 18'b000000001011100110; assign wn_im[116] = 18'b111111110100111111; 
assign wn_re[117] = 18'b000000001011100010; assign wn_im[117] = 18'b111111110100111010; 
assign wn_re[118] = 18'b000000001011011101; assign wn_im[118] = 18'b111111110100110101; 
assign wn_re[119] = 18'b000000001011011000; assign wn_im[119] = 18'b111111110100110000; 
assign wn_re[120] = 18'b000000001011010100; assign wn_im[120] = 18'b111111110100101011; 
assign wn_re[121] = 18'b000000001011001111; assign wn_im[121] = 18'b111111110100100111; 
assign wn_re[122] = 18'b000000001011001010; assign wn_im[122] = 18'b111111110100100010; 
assign wn_re[123] = 18'b000000001011000101; assign wn_im[123] = 18'b111111110100011101; 
assign wn_re[124] = 18'b000000001011000000; assign wn_im[124] = 18'b111111110100011001; 
assign wn_re[125] = 18'b000000001010111011; assign wn_im[125] = 18'b111111110100010100; 
assign wn_re[126] = 18'b000000001010110111; assign wn_im[126] = 18'b111111110100010000; 
assign wn_re[127] = 18'b000000001010110010; assign wn_im[127] = 18'b111111110100001011; 
assign wn_re[128] = 18'b000000001010101101; assign wn_im[128] = 18'b111111110100000111; 
assign wn_re[129] = 18'b000000001010101000; assign wn_im[129] = 18'b111111110100000010; 
assign wn_re[130] = 18'b000000001010100011; assign wn_im[130] = 18'b111111110011111110; 
assign wn_re[131] = 18'b000000001010011110; assign wn_im[131] = 18'b111111110011111001; 
assign wn_re[132] = 18'b000000001010011001; assign wn_im[132] = 18'b111111110011110101; 
assign wn_re[133] = 18'b000000001010010011; assign wn_im[133] = 18'b111111110011110001; 
assign wn_re[134] = 18'b000000001010001110; assign wn_im[134] = 18'b111111110011101100; 
assign wn_re[135] = 18'b000000001010001001; assign wn_im[135] = 18'b111111110011101000; 
assign wn_re[136] = 18'b000000001010000100; assign wn_im[136] = 18'b111111110011100100; 
assign wn_re[137] = 18'b000000001001111111; assign wn_im[137] = 18'b111111110011100000; 
assign wn_re[138] = 18'b000000001001111001; assign wn_im[138] = 18'b111111110011011011; 
assign wn_re[139] = 18'b000000001001110100; assign wn_im[139] = 18'b111111110011010111; 
assign wn_re[140] = 18'b000000001001101111; assign wn_im[140] = 18'b111111110011010011; 
assign wn_re[141] = 18'b000000001001101010; assign wn_im[141] = 18'b111111110011001111; 
assign wn_re[142] = 18'b000000001001100100; assign wn_im[142] = 18'b111111110011001011; 
assign wn_re[143] = 18'b000000001001011111; assign wn_im[143] = 18'b111111110011000111; 
assign wn_re[144] = 18'b000000001001011001; assign wn_im[144] = 18'b111111110011000011; 
assign wn_re[145] = 18'b000000001001010100; assign wn_im[145] = 18'b111111110010111111; 
assign wn_re[146] = 18'b000000001001001110; assign wn_im[146] = 18'b111111110010111011; 
assign wn_re[147] = 18'b000000001001001001; assign wn_im[147] = 18'b111111110010110111; 
assign wn_re[148] = 18'b000000001001000011; assign wn_im[148] = 18'b111111110010110100; 
assign wn_re[149] = 18'b000000001000111110; assign wn_im[149] = 18'b111111110010110000; 
assign wn_re[150] = 18'b000000001000111000; assign wn_im[150] = 18'b111111110010101100; 
assign wn_re[151] = 18'b000000001000110011; assign wn_im[151] = 18'b111111110010101000; 
assign wn_re[152] = 18'b000000001000101101; assign wn_im[152] = 18'b111111110010100101; 
assign wn_re[153] = 18'b000000001000101000; assign wn_im[153] = 18'b111111110010100001; 
assign wn_re[154] = 18'b000000001000100010; assign wn_im[154] = 18'b111111110010011101; 
assign wn_re[155] = 18'b000000001000011100; assign wn_im[155] = 18'b111111110010011010; 
assign wn_re[156] = 18'b000000001000010111; assign wn_im[156] = 18'b111111110010010110; 
assign wn_re[157] = 18'b000000001000010001; assign wn_im[157] = 18'b111111110010010011; 
assign wn_re[158] = 18'b000000001000001011; assign wn_im[158] = 18'b111111110010001111; 
assign wn_re[159] = 18'b000000001000000101; assign wn_im[159] = 18'b111111110010001100; 
assign wn_re[160] = 18'b000000001000000000; assign wn_im[160] = 18'b111111110010001001; 
assign wn_re[161] = 18'b000000000111111010; assign wn_im[161] = 18'b111111110010000101; 
assign wn_re[162] = 18'b000000000111110100; assign wn_im[162] = 18'b111111110010000010; 
assign wn_re[163] = 18'b000000000111101110; assign wn_im[163] = 18'b111111110001111111; 
assign wn_re[164] = 18'b000000000111101000; assign wn_im[164] = 18'b111111110001111100; 
assign wn_re[165] = 18'b000000000111100010; assign wn_im[165] = 18'b111111110001111000; 
assign wn_re[166] = 18'b000000000111011100; assign wn_im[166] = 18'b111111110001110101; 
assign wn_re[167] = 18'b000000000111010110; assign wn_im[167] = 18'b111111110001110010; 
assign wn_re[168] = 18'b000000000111010000; assign wn_im[168] = 18'b111111110001101111; 
assign wn_re[169] = 18'b000000000111001010; assign wn_im[169] = 18'b111111110001101100; 
assign wn_re[170] = 18'b000000000111000100; assign wn_im[170] = 18'b111111110001101001; 
assign wn_re[171] = 18'b000000000110111110; assign wn_im[171] = 18'b111111110001100110; 
assign wn_re[172] = 18'b000000000110111000; assign wn_im[172] = 18'b111111110001100011; 
assign wn_re[173] = 18'b000000000110110010; assign wn_im[173] = 18'b111111110001100000; 
assign wn_re[174] = 18'b000000000110101100; assign wn_im[174] = 18'b111111110001011110; 
assign wn_re[175] = 18'b000000000110100110; assign wn_im[175] = 18'b111111110001011011; 
assign wn_re[176] = 18'b000000000110100000; assign wn_im[176] = 18'b111111110001011000; 
assign wn_re[177] = 18'b000000000110011010; assign wn_im[177] = 18'b111111110001010101; 
assign wn_re[178] = 18'b000000000110010100; assign wn_im[178] = 18'b111111110001010011; 
assign wn_re[179] = 18'b000000000110001110; assign wn_im[179] = 18'b111111110001010000; 
assign wn_re[180] = 18'b000000000110000111; assign wn_im[180] = 18'b111111110001001101; 
assign wn_re[181] = 18'b000000000110000001; assign wn_im[181] = 18'b111111110001001011; 
assign wn_re[182] = 18'b000000000101111011; assign wn_im[182] = 18'b111111110001001000; 
assign wn_re[183] = 18'b000000000101110101; assign wn_im[183] = 18'b111111110001000110; 
assign wn_re[184] = 18'b000000000101101110; assign wn_im[184] = 18'b111111110001000100; 
assign wn_re[185] = 18'b000000000101101000; assign wn_im[185] = 18'b111111110001000001; 
assign wn_re[186] = 18'b000000000101100010; assign wn_im[186] = 18'b111111110000111111; 
assign wn_re[187] = 18'b000000000101011100; assign wn_im[187] = 18'b111111110000111100; 
assign wn_re[188] = 18'b000000000101010101; assign wn_im[188] = 18'b111111110000111010; 
assign wn_re[189] = 18'b000000000101001111; assign wn_im[189] = 18'b111111110000111000; 
assign wn_re[190] = 18'b000000000101001001; assign wn_im[190] = 18'b111111110000110110; 
assign wn_re[191] = 18'b000000000101000010; assign wn_im[191] = 18'b111111110000110100; 
assign wn_re[192] = 18'b000000000100111100; assign wn_im[192] = 18'b111111110000110010; 
assign wn_re[193] = 18'b000000000100110110; assign wn_im[193] = 18'b111111110000110000; 
assign wn_re[194] = 18'b000000000100101111; assign wn_im[194] = 18'b111111110000101110; 
assign wn_re[195] = 18'b000000000100101001; assign wn_im[195] = 18'b111111110000101100; 
assign wn_re[196] = 18'b000000000100100010; assign wn_im[196] = 18'b111111110000101010; 
assign wn_re[197] = 18'b000000000100011100; assign wn_im[197] = 18'b111111110000101000; 
assign wn_re[198] = 18'b000000000100010101; assign wn_im[198] = 18'b111111110000100110; 
assign wn_re[199] = 18'b000000000100001111; assign wn_im[199] = 18'b111111110000100100; 
assign wn_re[200] = 18'b000000000100001001; assign wn_im[200] = 18'b111111110000100010; 
assign wn_re[201] = 18'b000000000100000010; assign wn_im[201] = 18'b111111110000100001; 
assign wn_re[202] = 18'b000000000011111100; assign wn_im[202] = 18'b111111110000011111; 
assign wn_re[203] = 18'b000000000011110101; assign wn_im[203] = 18'b111111110000011101; 
assign wn_re[204] = 18'b000000000011101111; assign wn_im[204] = 18'b111111110000011100; 
assign wn_re[205] = 18'b000000000011101000; assign wn_im[205] = 18'b111111110000011010; 
assign wn_re[206] = 18'b000000000011100001; assign wn_im[206] = 18'b111111110000011001; 
assign wn_re[207] = 18'b000000000011011011; assign wn_im[207] = 18'b111111110000010111; 
assign wn_re[208] = 18'b000000000011010100; assign wn_im[208] = 18'b111111110000010110; 
assign wn_re[209] = 18'b000000000011001110; assign wn_im[209] = 18'b111111110000010101; 
assign wn_re[210] = 18'b000000000011000111; assign wn_im[210] = 18'b111111110000010011; 
assign wn_re[211] = 18'b000000000011000001; assign wn_im[211] = 18'b111111110000010010; 
assign wn_re[212] = 18'b000000000010111010; assign wn_im[212] = 18'b111111110000010001; 
assign wn_re[213] = 18'b000000000010110100; assign wn_im[213] = 18'b111111110000001111; 
assign wn_re[214] = 18'b000000000010101101; assign wn_im[214] = 18'b111111110000001110; 
assign wn_re[215] = 18'b000000000010100110; assign wn_im[215] = 18'b111111110000001101; 
assign wn_re[216] = 18'b000000000010100000; assign wn_im[216] = 18'b111111110000001100; 
assign wn_re[217] = 18'b000000000010011001; assign wn_im[217] = 18'b111111110000001011; 
assign wn_re[218] = 18'b000000000010010010; assign wn_im[218] = 18'b111111110000001010; 
assign wn_re[219] = 18'b000000000010001100; assign wn_im[219] = 18'b111111110000001001; 
assign wn_re[220] = 18'b000000000010000101; assign wn_im[220] = 18'b111111110000001000; 
assign wn_re[221] = 18'b000000000001111111; assign wn_im[221] = 18'b111111110000000111; 
assign wn_re[222] = 18'b000000000001111000; assign wn_im[222] = 18'b111111110000000111; 
assign wn_re[223] = 18'b000000000001110001; assign wn_im[223] = 18'b111111110000000110; 
assign wn_re[224] = 18'b000000000001101011; assign wn_im[224] = 18'b111111110000000101; 
assign wn_re[225] = 18'b000000000001100100; assign wn_im[225] = 18'b111111110000000100; 
assign wn_re[226] = 18'b000000000001011101; assign wn_im[226] = 18'b111111110000000100; 
assign wn_re[227] = 18'b000000000001010111; assign wn_im[227] = 18'b111111110000000011; 
assign wn_re[228] = 18'b000000000001010000; assign wn_im[228] = 18'b111111110000000011; 
assign wn_re[229] = 18'b000000000001001001; assign wn_im[229] = 18'b111111110000000010; 
assign wn_re[230] = 18'b000000000001000010; assign wn_im[230] = 18'b111111110000000010; 
assign wn_re[231] = 18'b000000000000111100; assign wn_im[231] = 18'b111111110000000001; 
assign wn_re[232] = 18'b000000000000110101; assign wn_im[232] = 18'b111111110000000001; 
assign wn_re[233] = 18'b000000000000101110; assign wn_im[233] = 18'b111111110000000001; 
assign wn_re[234] = 18'b000000000000101000; assign wn_im[234] = 18'b111111110000000000; 
assign wn_re[235] = 18'b000000000000100001; assign wn_im[235] = 18'b111111110000000000; 
assign wn_re[236] = 18'b000000000000011010; assign wn_im[236] = 18'b111111110000000000; 
assign wn_re[237] = 18'b000000000000010100; assign wn_im[237] = 18'b111111110000000000; 
assign wn_re[238] = 18'b000000000000001101; assign wn_im[238] = 18'b111111110000000000; 
assign wn_re[239] = 18'b000000000000000110; assign wn_im[239] = 18'b111111110000000000; 
assign wn_re[240] = 18'b000000000000000000; assign wn_im[240] = 18'b111111110000000000; 
assign wn_re[241] = 18'b111111111111111001; assign wn_im[241] = 18'b111111110000000000; 
assign wn_re[242] = 18'b111111111111110010; assign wn_im[242] = 18'b111111110000000000; 
assign wn_re[243] = 18'b111111111111101011; assign wn_im[243] = 18'b111111110000000000; 
assign wn_re[244] = 18'b111111111111100101; assign wn_im[244] = 18'b111111110000000000; 
assign wn_re[245] = 18'b111111111111011110; assign wn_im[245] = 18'b111111110000000000; 
assign wn_re[246] = 18'b111111111111010111; assign wn_im[246] = 18'b111111110000000000; 
assign wn_re[247] = 18'b111111111111010001; assign wn_im[247] = 18'b111111110000000001; 
assign wn_re[248] = 18'b111111111111001010; assign wn_im[248] = 18'b111111110000000001; 
assign wn_re[249] = 18'b111111111111000011; assign wn_im[249] = 18'b111111110000000001; 
assign wn_re[250] = 18'b111111111110111101; assign wn_im[250] = 18'b111111110000000010; 
assign wn_re[251] = 18'b111111111110110110; assign wn_im[251] = 18'b111111110000000010; 
assign wn_re[252] = 18'b111111111110101111; assign wn_im[252] = 18'b111111110000000011; 
assign wn_re[253] = 18'b111111111110101000; assign wn_im[253] = 18'b111111110000000011; 
assign wn_re[254] = 18'b111111111110100010; assign wn_im[254] = 18'b111111110000000100; 
assign wn_re[255] = 18'b111111111110011011; assign wn_im[255] = 18'b111111110000000100; 
assign wn_re[256] = 18'b111111111110010100; assign wn_im[256] = 18'b111111110000000101; 
assign wn_re[257] = 18'b111111111110001110; assign wn_im[257] = 18'b111111110000000110; 
assign wn_re[258] = 18'b111111111110000111; assign wn_im[258] = 18'b111111110000000111; 
assign wn_re[259] = 18'b111111111110000000; assign wn_im[259] = 18'b111111110000000111; 
assign wn_re[260] = 18'b111111111101111010; assign wn_im[260] = 18'b111111110000001000; 
assign wn_re[261] = 18'b111111111101110011; assign wn_im[261] = 18'b111111110000001001; 
assign wn_re[262] = 18'b111111111101101101; assign wn_im[262] = 18'b111111110000001010; 
assign wn_re[263] = 18'b111111111101100110; assign wn_im[263] = 18'b111111110000001011; 
assign wn_re[264] = 18'b111111111101011111; assign wn_im[264] = 18'b111111110000001100; 
assign wn_re[265] = 18'b111111111101011001; assign wn_im[265] = 18'b111111110000001101; 
assign wn_re[266] = 18'b111111111101010010; assign wn_im[266] = 18'b111111110000001110; 
assign wn_re[267] = 18'b111111111101001011; assign wn_im[267] = 18'b111111110000001111; 
assign wn_re[268] = 18'b111111111101000101; assign wn_im[268] = 18'b111111110000010001; 
assign wn_re[269] = 18'b111111111100111110; assign wn_im[269] = 18'b111111110000010010; 
assign wn_re[270] = 18'b111111111100111000; assign wn_im[270] = 18'b111111110000010011; 
assign wn_re[271] = 18'b111111111100110001; assign wn_im[271] = 18'b111111110000010101; 
assign wn_re[272] = 18'b111111111100101011; assign wn_im[272] = 18'b111111110000010110; 
assign wn_re[273] = 18'b111111111100100100; assign wn_im[273] = 18'b111111110000010111; 
assign wn_re[274] = 18'b111111111100011110; assign wn_im[274] = 18'b111111110000011001; 
assign wn_re[275] = 18'b111111111100010111; assign wn_im[275] = 18'b111111110000011010; 
assign wn_re[276] = 18'b111111111100010000; assign wn_im[276] = 18'b111111110000011100; 
assign wn_re[277] = 18'b111111111100001010; assign wn_im[277] = 18'b111111110000011101; 
assign wn_re[278] = 18'b111111111100000011; assign wn_im[278] = 18'b111111110000011111; 
assign wn_re[279] = 18'b111111111011111101; assign wn_im[279] = 18'b111111110000100001; 
assign wn_re[280] = 18'b111111111011110110; assign wn_im[280] = 18'b111111110000100010; 
assign wn_re[281] = 18'b111111111011110000; assign wn_im[281] = 18'b111111110000100100; 
assign wn_re[282] = 18'b111111111011101010; assign wn_im[282] = 18'b111111110000100110; 
assign wn_re[283] = 18'b111111111011100011; assign wn_im[283] = 18'b111111110000101000; 
assign wn_re[284] = 18'b111111111011011101; assign wn_im[284] = 18'b111111110000101010; 
assign wn_re[285] = 18'b111111111011010110; assign wn_im[285] = 18'b111111110000101100; 
assign wn_re[286] = 18'b111111111011010000; assign wn_im[286] = 18'b111111110000101110; 
assign wn_re[287] = 18'b111111111011001001; assign wn_im[287] = 18'b111111110000110000; 
assign wn_re[288] = 18'b111111111011000011; assign wn_im[288] = 18'b111111110000110010; 
assign wn_re[289] = 18'b111111111010111101; assign wn_im[289] = 18'b111111110000110100; 
assign wn_re[290] = 18'b111111111010110110; assign wn_im[290] = 18'b111111110000110110; 
assign wn_re[291] = 18'b111111111010110000; assign wn_im[291] = 18'b111111110000111000; 
assign wn_re[292] = 18'b111111111010101010; assign wn_im[292] = 18'b111111110000111010; 
assign wn_re[293] = 18'b111111111010100011; assign wn_im[293] = 18'b111111110000111100; 
assign wn_re[294] = 18'b111111111010011101; assign wn_im[294] = 18'b111111110000111111; 
assign wn_re[295] = 18'b111111111010010111; assign wn_im[295] = 18'b111111110001000001; 
assign wn_re[296] = 18'b111111111010010001; assign wn_im[296] = 18'b111111110001000100; 
assign wn_re[297] = 18'b111111111010001010; assign wn_im[297] = 18'b111111110001000110; 
assign wn_re[298] = 18'b111111111010000100; assign wn_im[298] = 18'b111111110001001000; 
assign wn_re[299] = 18'b111111111001111110; assign wn_im[299] = 18'b111111110001001011; 
assign wn_re[300] = 18'b111111111001111000; assign wn_im[300] = 18'b111111110001001101; 
assign wn_re[301] = 18'b111111111001110001; assign wn_im[301] = 18'b111111110001010000; 
assign wn_re[302] = 18'b111111111001101011; assign wn_im[302] = 18'b111111110001010011; 
assign wn_re[303] = 18'b111111111001100101; assign wn_im[303] = 18'b111111110001010101; 
assign wn_re[304] = 18'b111111111001011111; assign wn_im[304] = 18'b111111110001011000; 
assign wn_re[305] = 18'b111111111001011001; assign wn_im[305] = 18'b111111110001011011; 
assign wn_re[306] = 18'b111111111001010011; assign wn_im[306] = 18'b111111110001011110; 
assign wn_re[307] = 18'b111111111001001101; assign wn_im[307] = 18'b111111110001100000; 
assign wn_re[308] = 18'b111111111001000111; assign wn_im[308] = 18'b111111110001100011; 
assign wn_re[309] = 18'b111111111001000001; assign wn_im[309] = 18'b111111110001100110; 
assign wn_re[310] = 18'b111111111000111011; assign wn_im[310] = 18'b111111110001101001; 
assign wn_re[311] = 18'b111111111000110101; assign wn_im[311] = 18'b111111110001101100; 
assign wn_re[312] = 18'b111111111000101111; assign wn_im[312] = 18'b111111110001101111; 
assign wn_re[313] = 18'b111111111000101001; assign wn_im[313] = 18'b111111110001110010; 
assign wn_re[314] = 18'b111111111000100011; assign wn_im[314] = 18'b111111110001110101; 
assign wn_re[315] = 18'b111111111000011101; assign wn_im[315] = 18'b111111110001111000; 
assign wn_re[316] = 18'b111111111000010111; assign wn_im[316] = 18'b111111110001111100; 
assign wn_re[317] = 18'b111111111000010001; assign wn_im[317] = 18'b111111110001111111; 
assign wn_re[318] = 18'b111111111000001011; assign wn_im[318] = 18'b111111110010000010; 
assign wn_re[319] = 18'b111111111000000101; assign wn_im[319] = 18'b111111110010000101; 
assign wn_re[320] = 18'b111111111000000000; assign wn_im[320] = 18'b111111110010001001; 
assign wn_re[321] = 18'b111111110111111010; assign wn_im[321] = 18'b111111110010001100; 
assign wn_re[322] = 18'b111111110111110100; assign wn_im[322] = 18'b111111110010001111; 
assign wn_re[323] = 18'b111111110111101110; assign wn_im[323] = 18'b111111110010010011; 
assign wn_re[324] = 18'b111111110111101000; assign wn_im[324] = 18'b111111110010010110; 
assign wn_re[325] = 18'b111111110111100011; assign wn_im[325] = 18'b111111110010011010; 
assign wn_re[326] = 18'b111111110111011101; assign wn_im[326] = 18'b111111110010011101; 
assign wn_re[327] = 18'b111111110111010111; assign wn_im[327] = 18'b111111110010100001; 
assign wn_re[328] = 18'b111111110111010010; assign wn_im[328] = 18'b111111110010100101; 
assign wn_re[329] = 18'b111111110111001100; assign wn_im[329] = 18'b111111110010101000; 
assign wn_re[330] = 18'b111111110111000111; assign wn_im[330] = 18'b111111110010101100; 
assign wn_re[331] = 18'b111111110111000001; assign wn_im[331] = 18'b111111110010110000; 
assign wn_re[332] = 18'b111111110110111100; assign wn_im[332] = 18'b111111110010110100; 
assign wn_re[333] = 18'b111111110110110110; assign wn_im[333] = 18'b111111110010110111; 
assign wn_re[334] = 18'b111111110110110001; assign wn_im[334] = 18'b111111110010111011; 
assign wn_re[335] = 18'b111111110110101011; assign wn_im[335] = 18'b111111110010111111; 
assign wn_re[336] = 18'b111111110110100110; assign wn_im[336] = 18'b111111110011000011; 
assign wn_re[337] = 18'b111111110110100000; assign wn_im[337] = 18'b111111110011000111; 
assign wn_re[338] = 18'b111111110110011011; assign wn_im[338] = 18'b111111110011001011; 
assign wn_re[339] = 18'b111111110110010101; assign wn_im[339] = 18'b111111110011001111; 
assign wn_re[340] = 18'b111111110110010000; assign wn_im[340] = 18'b111111110011010011; 
assign wn_re[341] = 18'b111111110110001011; assign wn_im[341] = 18'b111111110011010111; 
assign wn_re[342] = 18'b111111110110000110; assign wn_im[342] = 18'b111111110011011011; 
assign wn_re[343] = 18'b111111110110000000; assign wn_im[343] = 18'b111111110011100000; 
assign wn_re[344] = 18'b111111110101111011; assign wn_im[344] = 18'b111111110011100100; 
assign wn_re[345] = 18'b111111110101110110; assign wn_im[345] = 18'b111111110011101000; 
assign wn_re[346] = 18'b111111110101110001; assign wn_im[346] = 18'b111111110011101100; 
assign wn_re[347] = 18'b111111110101101100; assign wn_im[347] = 18'b111111110011110001; 
assign wn_re[348] = 18'b111111110101100110; assign wn_im[348] = 18'b111111110011110101; 
assign wn_re[349] = 18'b111111110101100001; assign wn_im[349] = 18'b111111110011111001; 
assign wn_re[350] = 18'b111111110101011100; assign wn_im[350] = 18'b111111110011111110; 
assign wn_re[351] = 18'b111111110101010111; assign wn_im[351] = 18'b111111110100000010; 
assign wn_re[352] = 18'b111111110101010010; assign wn_im[352] = 18'b111111110100000111; 
assign wn_re[353] = 18'b111111110101001101; assign wn_im[353] = 18'b111111110100001011; 
assign wn_re[354] = 18'b111111110101001000; assign wn_im[354] = 18'b111111110100010000; 
assign wn_re[355] = 18'b111111110101000100; assign wn_im[355] = 18'b111111110100010100; 
assign wn_re[356] = 18'b111111110100111111; assign wn_im[356] = 18'b111111110100011001; 
assign wn_re[357] = 18'b111111110100111010; assign wn_im[357] = 18'b111111110100011101; 
assign wn_re[358] = 18'b111111110100110101; assign wn_im[358] = 18'b111111110100100010; 
assign wn_re[359] = 18'b111111110100110000; assign wn_im[359] = 18'b111111110100100111; 
assign wn_re[360] = 18'b111111110100101011; assign wn_im[360] = 18'b111111110100101011; 
assign wn_re[361] = 18'b111111110100100111; assign wn_im[361] = 18'b111111110100110000; 
assign wn_re[362] = 18'b111111110100100010; assign wn_im[362] = 18'b111111110100110101; 
assign wn_re[363] = 18'b111111110100011101; assign wn_im[363] = 18'b111111110100111010; 
assign wn_re[364] = 18'b111111110100011001; assign wn_im[364] = 18'b111111110100111111; 
assign wn_re[365] = 18'b111111110100010100; assign wn_im[365] = 18'b111111110101000100; 
assign wn_re[366] = 18'b111111110100010000; assign wn_im[366] = 18'b111111110101001000; 
assign wn_re[367] = 18'b111111110100001011; assign wn_im[367] = 18'b111111110101001101; 
assign wn_re[368] = 18'b111111110100000111; assign wn_im[368] = 18'b111111110101010010; 
assign wn_re[369] = 18'b111111110100000010; assign wn_im[369] = 18'b111111110101010111; 
assign wn_re[370] = 18'b111111110011111110; assign wn_im[370] = 18'b111111110101011100; 
assign wn_re[371] = 18'b111111110011111001; assign wn_im[371] = 18'b111111110101100001; 
assign wn_re[372] = 18'b111111110011110101; assign wn_im[372] = 18'b111111110101100110; 
assign wn_re[373] = 18'b111111110011110001; assign wn_im[373] = 18'b111111110101101100; 
assign wn_re[374] = 18'b111111110011101100; assign wn_im[374] = 18'b111111110101110001; 
assign wn_re[375] = 18'b111111110011101000; assign wn_im[375] = 18'b111111110101110110; 
assign wn_re[376] = 18'b111111110011100100; assign wn_im[376] = 18'b111111110101111011; 
assign wn_re[377] = 18'b111111110011100000; assign wn_im[377] = 18'b111111110110000000; 
assign wn_re[378] = 18'b111111110011011011; assign wn_im[378] = 18'b111111110110000110; 
assign wn_re[379] = 18'b111111110011010111; assign wn_im[379] = 18'b111111110110001011; 
assign wn_re[380] = 18'b111111110011010011; assign wn_im[380] = 18'b111111110110010000; 
assign wn_re[381] = 18'b111111110011001111; assign wn_im[381] = 18'b111111110110010101; 
assign wn_re[382] = 18'b111111110011001011; assign wn_im[382] = 18'b111111110110011011; 
assign wn_re[383] = 18'b111111110011000111; assign wn_im[383] = 18'b111111110110100000; 
assign wn_re[384] = 18'b111111110011000011; assign wn_im[384] = 18'b111111110110100110; 
assign wn_re[385] = 18'b111111110010111111; assign wn_im[385] = 18'b111111110110101011; 
assign wn_re[386] = 18'b111111110010111011; assign wn_im[386] = 18'b111111110110110001; 
assign wn_re[387] = 18'b111111110010110111; assign wn_im[387] = 18'b111111110110110110; 
assign wn_re[388] = 18'b111111110010110100; assign wn_im[388] = 18'b111111110110111100; 
assign wn_re[389] = 18'b111111110010110000; assign wn_im[389] = 18'b111111110111000001; 
assign wn_re[390] = 18'b111111110010101100; assign wn_im[390] = 18'b111111110111000111; 
assign wn_re[391] = 18'b111111110010101000; assign wn_im[391] = 18'b111111110111001100; 
assign wn_re[392] = 18'b111111110010100101; assign wn_im[392] = 18'b111111110111010010; 
assign wn_re[393] = 18'b111111110010100001; assign wn_im[393] = 18'b111111110111010111; 
assign wn_re[394] = 18'b111111110010011101; assign wn_im[394] = 18'b111111110111011101; 
assign wn_re[395] = 18'b111111110010011010; assign wn_im[395] = 18'b111111110111100011; 
assign wn_re[396] = 18'b111111110010010110; assign wn_im[396] = 18'b111111110111101000; 
assign wn_re[397] = 18'b111111110010010011; assign wn_im[397] = 18'b111111110111101110; 
assign wn_re[398] = 18'b111111110010001111; assign wn_im[398] = 18'b111111110111110100; 
assign wn_re[399] = 18'b111111110010001100; assign wn_im[399] = 18'b111111110111111010; 
assign wn_re[400] = 18'b111111110010001001; assign wn_im[400] = 18'b111111111000000000; 
assign wn_re[401] = 18'b111111110010000101; assign wn_im[401] = 18'b111111111000000101; 
assign wn_re[402] = 18'b111111110010000010; assign wn_im[402] = 18'b111111111000001011; 
assign wn_re[403] = 18'b111111110001111111; assign wn_im[403] = 18'b111111111000010001; 
assign wn_re[404] = 18'b111111110001111100; assign wn_im[404] = 18'b111111111000010111; 
assign wn_re[405] = 18'b111111110001111000; assign wn_im[405] = 18'b111111111000011101; 
assign wn_re[406] = 18'b111111110001110101; assign wn_im[406] = 18'b111111111000100011; 
assign wn_re[407] = 18'b111111110001110010; assign wn_im[407] = 18'b111111111000101001; 
assign wn_re[408] = 18'b111111110001101111; assign wn_im[408] = 18'b111111111000101111; 
assign wn_re[409] = 18'b111111110001101100; assign wn_im[409] = 18'b111111111000110101; 
assign wn_re[410] = 18'b111111110001101001; assign wn_im[410] = 18'b111111111000111011; 
assign wn_re[411] = 18'b111111110001100110; assign wn_im[411] = 18'b111111111001000001; 
assign wn_re[412] = 18'b111111110001100011; assign wn_im[412] = 18'b111111111001000111; 
assign wn_re[413] = 18'b111111110001100000; assign wn_im[413] = 18'b111111111001001101; 
assign wn_re[414] = 18'b111111110001011110; assign wn_im[414] = 18'b111111111001010011; 
assign wn_re[415] = 18'b111111110001011011; assign wn_im[415] = 18'b111111111001011001; 
assign wn_re[416] = 18'b111111110001011000; assign wn_im[416] = 18'b111111111001011111; 
assign wn_re[417] = 18'b111111110001010101; assign wn_im[417] = 18'b111111111001100101; 
assign wn_re[418] = 18'b111111110001010011; assign wn_im[418] = 18'b111111111001101011; 
assign wn_re[419] = 18'b111111110001010000; assign wn_im[419] = 18'b111111111001110001; 
assign wn_re[420] = 18'b111111110001001101; assign wn_im[420] = 18'b111111111001111000; 
assign wn_re[421] = 18'b111111110001001011; assign wn_im[421] = 18'b111111111001111110; 
assign wn_re[422] = 18'b111111110001001000; assign wn_im[422] = 18'b111111111010000100; 
assign wn_re[423] = 18'b111111110001000110; assign wn_im[423] = 18'b111111111010001010; 
assign wn_re[424] = 18'b111111110001000100; assign wn_im[424] = 18'b111111111010010001; 
assign wn_re[425] = 18'b111111110001000001; assign wn_im[425] = 18'b111111111010010111; 
assign wn_re[426] = 18'b111111110000111111; assign wn_im[426] = 18'b111111111010011101; 
assign wn_re[427] = 18'b111111110000111100; assign wn_im[427] = 18'b111111111010100011; 
assign wn_re[428] = 18'b111111110000111010; assign wn_im[428] = 18'b111111111010101010; 
assign wn_re[429] = 18'b111111110000111000; assign wn_im[429] = 18'b111111111010110000; 
assign wn_re[430] = 18'b111111110000110110; assign wn_im[430] = 18'b111111111010110110; 
assign wn_re[431] = 18'b111111110000110100; assign wn_im[431] = 18'b111111111010111101; 
assign wn_re[432] = 18'b111111110000110010; assign wn_im[432] = 18'b111111111011000011; 
assign wn_re[433] = 18'b111111110000110000; assign wn_im[433] = 18'b111111111011001001; 
assign wn_re[434] = 18'b111111110000101110; assign wn_im[434] = 18'b111111111011010000; 
assign wn_re[435] = 18'b111111110000101100; assign wn_im[435] = 18'b111111111011010110; 
assign wn_re[436] = 18'b111111110000101010; assign wn_im[436] = 18'b111111111011011101; 
assign wn_re[437] = 18'b111111110000101000; assign wn_im[437] = 18'b111111111011100011; 
assign wn_re[438] = 18'b111111110000100110; assign wn_im[438] = 18'b111111111011101010; 
assign wn_re[439] = 18'b111111110000100100; assign wn_im[439] = 18'b111111111011110000; 
assign wn_re[440] = 18'b111111110000100010; assign wn_im[440] = 18'b111111111011110110; 
assign wn_re[441] = 18'b111111110000100001; assign wn_im[441] = 18'b111111111011111101; 
assign wn_re[442] = 18'b111111110000011111; assign wn_im[442] = 18'b111111111100000011; 
assign wn_re[443] = 18'b111111110000011101; assign wn_im[443] = 18'b111111111100001010; 
assign wn_re[444] = 18'b111111110000011100; assign wn_im[444] = 18'b111111111100010000; 
assign wn_re[445] = 18'b111111110000011010; assign wn_im[445] = 18'b111111111100010111; 
assign wn_re[446] = 18'b111111110000011001; assign wn_im[446] = 18'b111111111100011110; 
assign wn_re[447] = 18'b111111110000010111; assign wn_im[447] = 18'b111111111100100100; 
assign wn_re[448] = 18'b111111110000010110; assign wn_im[448] = 18'b111111111100101011; 
assign wn_re[449] = 18'b111111110000010101; assign wn_im[449] = 18'b111111111100110001; 
assign wn_re[450] = 18'b111111110000010011; assign wn_im[450] = 18'b111111111100111000; 
assign wn_re[451] = 18'b111111110000010010; assign wn_im[451] = 18'b111111111100111110; 
assign wn_re[452] = 18'b111111110000010001; assign wn_im[452] = 18'b111111111101000101; 
assign wn_re[453] = 18'b111111110000001111; assign wn_im[453] = 18'b111111111101001011; 
assign wn_re[454] = 18'b111111110000001110; assign wn_im[454] = 18'b111111111101010010; 
assign wn_re[455] = 18'b111111110000001101; assign wn_im[455] = 18'b111111111101011001; 
assign wn_re[456] = 18'b111111110000001100; assign wn_im[456] = 18'b111111111101011111; 
assign wn_re[457] = 18'b111111110000001011; assign wn_im[457] = 18'b111111111101100110; 
assign wn_re[458] = 18'b111111110000001010; assign wn_im[458] = 18'b111111111101101101; 
assign wn_re[459] = 18'b111111110000001001; assign wn_im[459] = 18'b111111111101110011; 
assign wn_re[460] = 18'b111111110000001000; assign wn_im[460] = 18'b111111111101111010; 
assign wn_re[461] = 18'b111111110000000111; assign wn_im[461] = 18'b111111111110000000; 
assign wn_re[462] = 18'b111111110000000111; assign wn_im[462] = 18'b111111111110000111; 
assign wn_re[463] = 18'b111111110000000110; assign wn_im[463] = 18'b111111111110001110; 
assign wn_re[464] = 18'b111111110000000101; assign wn_im[464] = 18'b111111111110010100; 
assign wn_re[465] = 18'b111111110000000100; assign wn_im[465] = 18'b111111111110011011; 
assign wn_re[466] = 18'b111111110000000100; assign wn_im[466] = 18'b111111111110100010; 
assign wn_re[467] = 18'b111111110000000011; assign wn_im[467] = 18'b111111111110101000; 
assign wn_re[468] = 18'b111111110000000011; assign wn_im[468] = 18'b111111111110101111; 
assign wn_re[469] = 18'b111111110000000010; assign wn_im[469] = 18'b111111111110110110; 
assign wn_re[470] = 18'b111111110000000010; assign wn_im[470] = 18'b111111111110111101; 
assign wn_re[471] = 18'b111111110000000001; assign wn_im[471] = 18'b111111111111000011; 
assign wn_re[472] = 18'b111111110000000001; assign wn_im[472] = 18'b111111111111001010; 
assign wn_re[473] = 18'b111111110000000001; assign wn_im[473] = 18'b111111111111010001; 
assign wn_re[474] = 18'b111111110000000000; assign wn_im[474] = 18'b111111111111010111; 
assign wn_re[475] = 18'b111111110000000000; assign wn_im[475] = 18'b111111111111011110; 
assign wn_re[476] = 18'b111111110000000000; assign wn_im[476] = 18'b111111111111100101; 
assign wn_re[477] = 18'b111111110000000000; assign wn_im[477] = 18'b111111111111101011; 
assign wn_re[478] = 18'b111111110000000000; assign wn_im[478] = 18'b111111111111110010; 
assign wn_re[479] = 18'b111111110000000000; assign wn_im[479] = 18'b111111111111111001; 
assign wn_re[480] = 18'b111111110000000000; assign wn_im[480] = 18'b111111111111111111; 
assign wn_re[481] = 18'b111111110000000000; assign wn_im[481] = 18'b000000000000000110; 
assign wn_re[482] = 18'b111111110000000000; assign wn_im[482] = 18'b000000000000001101; 
assign wn_re[483] = 18'b111111110000000000; assign wn_im[483] = 18'b000000000000010100; 
assign wn_re[484] = 18'b111111110000000000; assign wn_im[484] = 18'b000000000000011010; 
assign wn_re[485] = 18'b111111110000000000; assign wn_im[485] = 18'b000000000000100001; 
assign wn_re[486] = 18'b111111110000000000; assign wn_im[486] = 18'b000000000000101000; 
assign wn_re[487] = 18'b111111110000000001; assign wn_im[487] = 18'b000000000000101110; 
assign wn_re[488] = 18'b111111110000000001; assign wn_im[488] = 18'b000000000000110101; 
assign wn_re[489] = 18'b111111110000000001; assign wn_im[489] = 18'b000000000000111100; 
assign wn_re[490] = 18'b111111110000000010; assign wn_im[490] = 18'b000000000001000010; 
assign wn_re[491] = 18'b111111110000000010; assign wn_im[491] = 18'b000000000001001001; 
assign wn_re[492] = 18'b111111110000000011; assign wn_im[492] = 18'b000000000001010000; 
assign wn_re[493] = 18'b111111110000000011; assign wn_im[493] = 18'b000000000001010111; 
assign wn_re[494] = 18'b111111110000000100; assign wn_im[494] = 18'b000000000001011101; 
assign wn_re[495] = 18'b111111110000000100; assign wn_im[495] = 18'b000000000001100100; 
assign wn_re[496] = 18'b111111110000000101; assign wn_im[496] = 18'b000000000001101011; 
assign wn_re[497] = 18'b111111110000000110; assign wn_im[497] = 18'b000000000001110001; 
assign wn_re[498] = 18'b111111110000000111; assign wn_im[498] = 18'b000000000001111000; 
assign wn_re[499] = 18'b111111110000000111; assign wn_im[499] = 18'b000000000001111111; 
assign wn_re[500] = 18'b111111110000001000; assign wn_im[500] = 18'b000000000010000101; 
assign wn_re[501] = 18'b111111110000001001; assign wn_im[501] = 18'b000000000010001100; 
assign wn_re[502] = 18'b111111110000001010; assign wn_im[502] = 18'b000000000010010010; 
assign wn_re[503] = 18'b111111110000001011; assign wn_im[503] = 18'b000000000010011001; 
assign wn_re[504] = 18'b111111110000001100; assign wn_im[504] = 18'b000000000010100000; 
assign wn_re[505] = 18'b111111110000001101; assign wn_im[505] = 18'b000000000010100110; 
assign wn_re[506] = 18'b111111110000001110; assign wn_im[506] = 18'b000000000010101101; 
assign wn_re[507] = 18'b111111110000001111; assign wn_im[507] = 18'b000000000010110100; 
assign wn_re[508] = 18'b111111110000010001; assign wn_im[508] = 18'b000000000010111010; 
assign wn_re[509] = 18'b111111110000010010; assign wn_im[509] = 18'b000000000011000001; 
assign wn_re[510] = 18'b111111110000010011; assign wn_im[510] = 18'b000000000011000111; 
assign wn_re[511] = 18'b111111110000010101; assign wn_im[511] = 18'b000000000011001110; 
assign wn_re[512] = 18'b111111110000010110; assign wn_im[512] = 18'b000000000011010100; 
assign wn_re[513] = 18'b111111110000010111; assign wn_im[513] = 18'b000000000011011011; 
assign wn_re[514] = 18'b111111110000011001; assign wn_im[514] = 18'b000000000011100001; 
assign wn_re[515] = 18'b111111110000011010; assign wn_im[515] = 18'b000000000011101000; 
assign wn_re[516] = 18'b111111110000011100; assign wn_im[516] = 18'b000000000011101111; 
assign wn_re[517] = 18'b111111110000011101; assign wn_im[517] = 18'b000000000011110101; 
assign wn_re[518] = 18'b111111110000011111; assign wn_im[518] = 18'b000000000011111100; 
assign wn_re[519] = 18'b111111110000100001; assign wn_im[519] = 18'b000000000100000010; 
assign wn_re[520] = 18'b111111110000100010; assign wn_im[520] = 18'b000000000100001001; 
assign wn_re[521] = 18'b111111110000100100; assign wn_im[521] = 18'b000000000100001111; 
assign wn_re[522] = 18'b111111110000100110; assign wn_im[522] = 18'b000000000100010101; 
assign wn_re[523] = 18'b111111110000101000; assign wn_im[523] = 18'b000000000100011100; 
assign wn_re[524] = 18'b111111110000101010; assign wn_im[524] = 18'b000000000100100010; 
assign wn_re[525] = 18'b111111110000101100; assign wn_im[525] = 18'b000000000100101001; 
assign wn_re[526] = 18'b111111110000101110; assign wn_im[526] = 18'b000000000100101111; 
assign wn_re[527] = 18'b111111110000110000; assign wn_im[527] = 18'b000000000100110110; 
assign wn_re[528] = 18'b111111110000110010; assign wn_im[528] = 18'b000000000100111100; 
assign wn_re[529] = 18'b111111110000110100; assign wn_im[529] = 18'b000000000101000010; 
assign wn_re[530] = 18'b111111110000110110; assign wn_im[530] = 18'b000000000101001001; 
assign wn_re[531] = 18'b111111110000111000; assign wn_im[531] = 18'b000000000101001111; 
assign wn_re[532] = 18'b111111110000111010; assign wn_im[532] = 18'b000000000101010101; 
assign wn_re[533] = 18'b111111110000111100; assign wn_im[533] = 18'b000000000101011100; 
assign wn_re[534] = 18'b111111110000111111; assign wn_im[534] = 18'b000000000101100010; 
assign wn_re[535] = 18'b111111110001000001; assign wn_im[535] = 18'b000000000101101000; 
assign wn_re[536] = 18'b111111110001000100; assign wn_im[536] = 18'b000000000101101110; 
assign wn_re[537] = 18'b111111110001000110; assign wn_im[537] = 18'b000000000101110101; 
assign wn_re[538] = 18'b111111110001001000; assign wn_im[538] = 18'b000000000101111011; 
assign wn_re[539] = 18'b111111110001001011; assign wn_im[539] = 18'b000000000110000001; 
assign wn_re[540] = 18'b111111110001001101; assign wn_im[540] = 18'b000000000110000111; 
assign wn_re[541] = 18'b111111110001010000; assign wn_im[541] = 18'b000000000110001110; 
assign wn_re[542] = 18'b111111110001010011; assign wn_im[542] = 18'b000000000110010100; 
assign wn_re[543] = 18'b111111110001010101; assign wn_im[543] = 18'b000000000110011010; 
assign wn_re[544] = 18'b111111110001011000; assign wn_im[544] = 18'b000000000110100000; 
assign wn_re[545] = 18'b111111110001011011; assign wn_im[545] = 18'b000000000110100110; 
assign wn_re[546] = 18'b111111110001011110; assign wn_im[546] = 18'b000000000110101100; 
assign wn_re[547] = 18'b111111110001100000; assign wn_im[547] = 18'b000000000110110010; 
assign wn_re[548] = 18'b111111110001100011; assign wn_im[548] = 18'b000000000110111000; 
assign wn_re[549] = 18'b111111110001100110; assign wn_im[549] = 18'b000000000110111110; 
assign wn_re[550] = 18'b111111110001101001; assign wn_im[550] = 18'b000000000111000100; 
assign wn_re[551] = 18'b111111110001101100; assign wn_im[551] = 18'b000000000111001010; 
assign wn_re[552] = 18'b111111110001101111; assign wn_im[552] = 18'b000000000111010000; 
assign wn_re[553] = 18'b111111110001110010; assign wn_im[553] = 18'b000000000111010110; 
assign wn_re[554] = 18'b111111110001110101; assign wn_im[554] = 18'b000000000111011100; 
assign wn_re[555] = 18'b111111110001111000; assign wn_im[555] = 18'b000000000111100010; 
assign wn_re[556] = 18'b111111110001111100; assign wn_im[556] = 18'b000000000111101000; 
assign wn_re[557] = 18'b111111110001111111; assign wn_im[557] = 18'b000000000111101110; 
assign wn_re[558] = 18'b111111110010000010; assign wn_im[558] = 18'b000000000111110100; 
assign wn_re[559] = 18'b111111110010000101; assign wn_im[559] = 18'b000000000111111010; 
assign wn_re[560] = 18'b111111110010001001; assign wn_im[560] = 18'b000000000111111111; 
assign wn_re[561] = 18'b111111110010001100; assign wn_im[561] = 18'b000000001000000101; 
assign wn_re[562] = 18'b111111110010001111; assign wn_im[562] = 18'b000000001000001011; 
assign wn_re[563] = 18'b111111110010010011; assign wn_im[563] = 18'b000000001000010001; 
assign wn_re[564] = 18'b111111110010010110; assign wn_im[564] = 18'b000000001000010111; 
assign wn_re[565] = 18'b111111110010011010; assign wn_im[565] = 18'b000000001000011100; 
assign wn_re[566] = 18'b111111110010011101; assign wn_im[566] = 18'b000000001000100010; 
assign wn_re[567] = 18'b111111110010100001; assign wn_im[567] = 18'b000000001000101000; 
assign wn_re[568] = 18'b111111110010100101; assign wn_im[568] = 18'b000000001000101101; 
assign wn_re[569] = 18'b111111110010101000; assign wn_im[569] = 18'b000000001000110011; 
assign wn_re[570] = 18'b111111110010101100; assign wn_im[570] = 18'b000000001000111000; 
assign wn_re[571] = 18'b111111110010110000; assign wn_im[571] = 18'b000000001000111110; 
assign wn_re[572] = 18'b111111110010110100; assign wn_im[572] = 18'b000000001001000011; 
assign wn_re[573] = 18'b111111110010110111; assign wn_im[573] = 18'b000000001001001001; 
assign wn_re[574] = 18'b111111110010111011; assign wn_im[574] = 18'b000000001001001110; 
assign wn_re[575] = 18'b111111110010111111; assign wn_im[575] = 18'b000000001001010100; 
assign wn_re[576] = 18'b111111110011000011; assign wn_im[576] = 18'b000000001001011001; 
assign wn_re[577] = 18'b111111110011000111; assign wn_im[577] = 18'b000000001001011111; 
assign wn_re[578] = 18'b111111110011001011; assign wn_im[578] = 18'b000000001001100100; 
assign wn_re[579] = 18'b111111110011001111; assign wn_im[579] = 18'b000000001001101010; 
assign wn_re[580] = 18'b111111110011010011; assign wn_im[580] = 18'b000000001001101111; 
assign wn_re[581] = 18'b111111110011010111; assign wn_im[581] = 18'b000000001001110100; 
assign wn_re[582] = 18'b111111110011011011; assign wn_im[582] = 18'b000000001001111001; 
assign wn_re[583] = 18'b111111110011100000; assign wn_im[583] = 18'b000000001001111111; 
assign wn_re[584] = 18'b111111110011100100; assign wn_im[584] = 18'b000000001010000100; 
assign wn_re[585] = 18'b111111110011101000; assign wn_im[585] = 18'b000000001010001001; 
assign wn_re[586] = 18'b111111110011101100; assign wn_im[586] = 18'b000000001010001110; 
assign wn_re[587] = 18'b111111110011110001; assign wn_im[587] = 18'b000000001010010011; 
assign wn_re[588] = 18'b111111110011110101; assign wn_im[588] = 18'b000000001010011001; 
assign wn_re[589] = 18'b111111110011111001; assign wn_im[589] = 18'b000000001010011110; 
assign wn_re[590] = 18'b111111110011111110; assign wn_im[590] = 18'b000000001010100011; 
assign wn_re[591] = 18'b111111110100000010; assign wn_im[591] = 18'b000000001010101000; 
assign wn_re[592] = 18'b111111110100000111; assign wn_im[592] = 18'b000000001010101101; 
assign wn_re[593] = 18'b111111110100001011; assign wn_im[593] = 18'b000000001010110010; 
assign wn_re[594] = 18'b111111110100010000; assign wn_im[594] = 18'b000000001010110111; 
assign wn_re[595] = 18'b111111110100010100; assign wn_im[595] = 18'b000000001010111011; 
assign wn_re[596] = 18'b111111110100011001; assign wn_im[596] = 18'b000000001011000000; 
assign wn_re[597] = 18'b111111110100011101; assign wn_im[597] = 18'b000000001011000101; 
assign wn_re[598] = 18'b111111110100100010; assign wn_im[598] = 18'b000000001011001010; 
assign wn_re[599] = 18'b111111110100100111; assign wn_im[599] = 18'b000000001011001111; 
assign wn_re[600] = 18'b111111110100101011; assign wn_im[600] = 18'b000000001011010100; 
assign wn_re[601] = 18'b111111110100110000; assign wn_im[601] = 18'b000000001011011000; 
assign wn_re[602] = 18'b111111110100110101; assign wn_im[602] = 18'b000000001011011101; 
assign wn_re[603] = 18'b111111110100111010; assign wn_im[603] = 18'b000000001011100010; 
assign wn_re[604] = 18'b111111110100111111; assign wn_im[604] = 18'b000000001011100110; 
assign wn_re[605] = 18'b111111110101000100; assign wn_im[605] = 18'b000000001011101011; 
assign wn_re[606] = 18'b111111110101001000; assign wn_im[606] = 18'b000000001011101111; 
assign wn_re[607] = 18'b111111110101001101; assign wn_im[607] = 18'b000000001011110100; 
assign wn_re[608] = 18'b111111110101010010; assign wn_im[608] = 18'b000000001011111000; 
assign wn_re[609] = 18'b111111110101010111; assign wn_im[609] = 18'b000000001011111101; 
assign wn_re[610] = 18'b111111110101011100; assign wn_im[610] = 18'b000000001100000001; 
assign wn_re[611] = 18'b111111110101100001; assign wn_im[611] = 18'b000000001100000110; 
assign wn_re[612] = 18'b111111110101100110; assign wn_im[612] = 18'b000000001100001010; 
assign wn_re[613] = 18'b111111110101101100; assign wn_im[613] = 18'b000000001100001110; 
assign wn_re[614] = 18'b111111110101110001; assign wn_im[614] = 18'b000000001100010011; 
assign wn_re[615] = 18'b111111110101110110; assign wn_im[615] = 18'b000000001100010111; 
assign wn_re[616] = 18'b111111110101111011; assign wn_im[616] = 18'b000000001100011011; 
assign wn_re[617] = 18'b111111110110000000; assign wn_im[617] = 18'b000000001100011111; 
assign wn_re[618] = 18'b111111110110000110; assign wn_im[618] = 18'b000000001100100100; 
assign wn_re[619] = 18'b111111110110001011; assign wn_im[619] = 18'b000000001100101000; 
assign wn_re[620] = 18'b111111110110010000; assign wn_im[620] = 18'b000000001100101100; 
assign wn_re[621] = 18'b111111110110010101; assign wn_im[621] = 18'b000000001100110000; 
assign wn_re[622] = 18'b111111110110011011; assign wn_im[622] = 18'b000000001100110100; 
assign wn_re[623] = 18'b111111110110100000; assign wn_im[623] = 18'b000000001100111000; 
assign wn_re[624] = 18'b111111110110100110; assign wn_im[624] = 18'b000000001100111100; 
assign wn_re[625] = 18'b111111110110101011; assign wn_im[625] = 18'b000000001101000000; 
assign wn_re[626] = 18'b111111110110110001; assign wn_im[626] = 18'b000000001101000100; 
assign wn_re[627] = 18'b111111110110110110; assign wn_im[627] = 18'b000000001101001000; 
assign wn_re[628] = 18'b111111110110111100; assign wn_im[628] = 18'b000000001101001011; 
assign wn_re[629] = 18'b111111110111000001; assign wn_im[629] = 18'b000000001101001111; 
assign wn_re[630] = 18'b111111110111000111; assign wn_im[630] = 18'b000000001101010011; 
assign wn_re[631] = 18'b111111110111001100; assign wn_im[631] = 18'b000000001101010111; 
assign wn_re[632] = 18'b111111110111010010; assign wn_im[632] = 18'b000000001101011010; 
assign wn_re[633] = 18'b111111110111010111; assign wn_im[633] = 18'b000000001101011110; 
assign wn_re[634] = 18'b111111110111011101; assign wn_im[634] = 18'b000000001101100010; 
assign wn_re[635] = 18'b111111110111100011; assign wn_im[635] = 18'b000000001101100101; 
assign wn_re[636] = 18'b111111110111101000; assign wn_im[636] = 18'b000000001101101001; 
assign wn_re[637] = 18'b111111110111101110; assign wn_im[637] = 18'b000000001101101100; 
assign wn_re[638] = 18'b111111110111110100; assign wn_im[638] = 18'b000000001101110000; 
assign wn_re[639] = 18'b111111110111111010; assign wn_im[639] = 18'b000000001101110011; 
assign wn_re[640] = 18'b111111110111111111; assign wn_im[640] = 18'b000000001101110110; 
assign wn_re[641] = 18'b111111111000000101; assign wn_im[641] = 18'b000000001101111010; 
assign wn_re[642] = 18'b111111111000001011; assign wn_im[642] = 18'b000000001101111101; 
assign wn_re[643] = 18'b111111111000010001; assign wn_im[643] = 18'b000000001110000000; 
assign wn_re[644] = 18'b111111111000010111; assign wn_im[644] = 18'b000000001110000011; 
assign wn_re[645] = 18'b111111111000011101; assign wn_im[645] = 18'b000000001110000111; 
assign wn_re[646] = 18'b111111111000100011; assign wn_im[646] = 18'b000000001110001010; 
assign wn_re[647] = 18'b111111111000101001; assign wn_im[647] = 18'b000000001110001101; 
assign wn_re[648] = 18'b111111111000101111; assign wn_im[648] = 18'b000000001110010000; 
assign wn_re[649] = 18'b111111111000110101; assign wn_im[649] = 18'b000000001110010011; 
assign wn_re[650] = 18'b111111111000111011; assign wn_im[650] = 18'b000000001110010110; 
assign wn_re[651] = 18'b111111111001000001; assign wn_im[651] = 18'b000000001110011001; 
assign wn_re[652] = 18'b111111111001000111; assign wn_im[652] = 18'b000000001110011100; 
assign wn_re[653] = 18'b111111111001001101; assign wn_im[653] = 18'b000000001110011111; 
assign wn_re[654] = 18'b111111111001010011; assign wn_im[654] = 18'b000000001110100001; 
assign wn_re[655] = 18'b111111111001011001; assign wn_im[655] = 18'b000000001110100100; 
assign wn_re[656] = 18'b111111111001011111; assign wn_im[656] = 18'b000000001110100111; 
assign wn_re[657] = 18'b111111111001100101; assign wn_im[657] = 18'b000000001110101010; 
assign wn_re[658] = 18'b111111111001101011; assign wn_im[658] = 18'b000000001110101100; 
assign wn_re[659] = 18'b111111111001110001; assign wn_im[659] = 18'b000000001110101111; 
assign wn_re[660] = 18'b111111111001111000; assign wn_im[660] = 18'b000000001110110010; 
assign wn_re[661] = 18'b111111111001111110; assign wn_im[661] = 18'b000000001110110100; 
assign wn_re[662] = 18'b111111111010000100; assign wn_im[662] = 18'b000000001110110111; 
assign wn_re[663] = 18'b111111111010001010; assign wn_im[663] = 18'b000000001110111001; 
assign wn_re[664] = 18'b111111111010010001; assign wn_im[664] = 18'b000000001110111011; 
assign wn_re[665] = 18'b111111111010010111; assign wn_im[665] = 18'b000000001110111110; 
assign wn_re[666] = 18'b111111111010011101; assign wn_im[666] = 18'b000000001111000000; 
assign wn_re[667] = 18'b111111111010100011; assign wn_im[667] = 18'b000000001111000011; 
assign wn_re[668] = 18'b111111111010101010; assign wn_im[668] = 18'b000000001111000101; 
assign wn_re[669] = 18'b111111111010110000; assign wn_im[669] = 18'b000000001111000111; 
assign wn_re[670] = 18'b111111111010110110; assign wn_im[670] = 18'b000000001111001001; 
assign wn_re[671] = 18'b111111111010111101; assign wn_im[671] = 18'b000000001111001011; 
assign wn_re[672] = 18'b111111111011000011; assign wn_im[672] = 18'b000000001111001101; 
assign wn_re[673] = 18'b111111111011001001; assign wn_im[673] = 18'b000000001111001111; 
assign wn_re[674] = 18'b111111111011010000; assign wn_im[674] = 18'b000000001111010001; 
assign wn_re[675] = 18'b111111111011010110; assign wn_im[675] = 18'b000000001111010011; 
assign wn_re[676] = 18'b111111111011011101; assign wn_im[676] = 18'b000000001111010101; 
assign wn_re[677] = 18'b111111111011100011; assign wn_im[677] = 18'b000000001111010111; 
assign wn_re[678] = 18'b111111111011101010; assign wn_im[678] = 18'b000000001111011001; 
assign wn_re[679] = 18'b111111111011110000; assign wn_im[679] = 18'b000000001111011011; 
assign wn_re[680] = 18'b111111111011110110; assign wn_im[680] = 18'b000000001111011101; 
assign wn_re[681] = 18'b111111111011111101; assign wn_im[681] = 18'b000000001111011110; 
assign wn_re[682] = 18'b111111111100000011; assign wn_im[682] = 18'b000000001111100000; 
assign wn_re[683] = 18'b111111111100001010; assign wn_im[683] = 18'b000000001111100010; 
assign wn_re[684] = 18'b111111111100010000; assign wn_im[684] = 18'b000000001111100011; 
assign wn_re[685] = 18'b111111111100010111; assign wn_im[685] = 18'b000000001111100101; 
assign wn_re[686] = 18'b111111111100011110; assign wn_im[686] = 18'b000000001111100110; 
assign wn_re[687] = 18'b111111111100100100; assign wn_im[687] = 18'b000000001111101000; 
assign wn_re[688] = 18'b111111111100101011; assign wn_im[688] = 18'b000000001111101001; 
assign wn_re[689] = 18'b111111111100110001; assign wn_im[689] = 18'b000000001111101010; 
assign wn_re[690] = 18'b111111111100111000; assign wn_im[690] = 18'b000000001111101100; 
assign wn_re[691] = 18'b111111111100111110; assign wn_im[691] = 18'b000000001111101101; 
assign wn_re[692] = 18'b111111111101000101; assign wn_im[692] = 18'b000000001111101110; 
assign wn_re[693] = 18'b111111111101001011; assign wn_im[693] = 18'b000000001111110000; 
assign wn_re[694] = 18'b111111111101010010; assign wn_im[694] = 18'b000000001111110001; 
assign wn_re[695] = 18'b111111111101011001; assign wn_im[695] = 18'b000000001111110010; 
assign wn_re[696] = 18'b111111111101011111; assign wn_im[696] = 18'b000000001111110011; 
assign wn_re[697] = 18'b111111111101100110; assign wn_im[697] = 18'b000000001111110100; 
assign wn_re[698] = 18'b111111111101101101; assign wn_im[698] = 18'b000000001111110101; 
assign wn_re[699] = 18'b111111111101110011; assign wn_im[699] = 18'b000000001111110110; 
assign wn_re[700] = 18'b111111111101111010; assign wn_im[700] = 18'b000000001111110111; 
assign wn_re[701] = 18'b111111111110000000; assign wn_im[701] = 18'b000000001111111000; 
assign wn_re[702] = 18'b111111111110000111; assign wn_im[702] = 18'b000000001111111000; 
assign wn_re[703] = 18'b111111111110001110; assign wn_im[703] = 18'b000000001111111001; 
assign wn_re[704] = 18'b111111111110010100; assign wn_im[704] = 18'b000000001111111010; 
assign wn_re[705] = 18'b111111111110011011; assign wn_im[705] = 18'b000000001111111011; 
assign wn_re[706] = 18'b111111111110100010; assign wn_im[706] = 18'b000000001111111011; 
assign wn_re[707] = 18'b111111111110101000; assign wn_im[707] = 18'b000000001111111100; 
assign wn_re[708] = 18'b111111111110101111; assign wn_im[708] = 18'b000000001111111100; 
assign wn_re[709] = 18'b111111111110110110; assign wn_im[709] = 18'b000000001111111101; 
assign wn_re[710] = 18'b111111111110111101; assign wn_im[710] = 18'b000000001111111101; 
assign wn_re[711] = 18'b111111111111000011; assign wn_im[711] = 18'b000000001111111110; 
assign wn_re[712] = 18'b111111111111001010; assign wn_im[712] = 18'b000000001111111110; 
assign wn_re[713] = 18'b111111111111010001; assign wn_im[713] = 18'b000000001111111110; 
assign wn_re[714] = 18'b111111111111010111; assign wn_im[714] = 18'b000000001111111111; 
assign wn_re[715] = 18'b111111111111011110; assign wn_im[715] = 18'b000000001111111111; 
assign wn_re[716] = 18'b111111111111100101; assign wn_im[716] = 18'b000000001111111111; 
assign wn_re[717] = 18'b111111111111101011; assign wn_im[717] = 18'b000000001111111111; 
assign wn_re[718] = 18'b111111111111110010; assign wn_im[718] = 18'b000000001111111111; 
assign wn_re[719] = 18'b111111111111111001; assign wn_im[719] = 18'b000000001111111111; 
assign wn_re[720] = 18'b111111111111111111; assign wn_im[720] = 18'b000000010000000000; 
assign wn_re[721] = 18'b000000000000000110; assign wn_im[721] = 18'b000000001111111111; 
assign wn_re[722] = 18'b000000000000001101; assign wn_im[722] = 18'b000000001111111111; 
assign wn_re[723] = 18'b000000000000010100; assign wn_im[723] = 18'b000000001111111111; 
assign wn_re[724] = 18'b000000000000011010; assign wn_im[724] = 18'b000000001111111111; 
assign wn_re[725] = 18'b000000000000100001; assign wn_im[725] = 18'b000000001111111111; 
assign wn_re[726] = 18'b000000000000101000; assign wn_im[726] = 18'b000000001111111111; 
assign wn_re[727] = 18'b000000000000101110; assign wn_im[727] = 18'b000000001111111110; 
assign wn_re[728] = 18'b000000000000110101; assign wn_im[728] = 18'b000000001111111110; 
assign wn_re[729] = 18'b000000000000111100; assign wn_im[729] = 18'b000000001111111110; 
assign wn_re[730] = 18'b000000000001000010; assign wn_im[730] = 18'b000000001111111101; 
assign wn_re[731] = 18'b000000000001001001; assign wn_im[731] = 18'b000000001111111101; 
assign wn_re[732] = 18'b000000000001010000; assign wn_im[732] = 18'b000000001111111100; 
assign wn_re[733] = 18'b000000000001010111; assign wn_im[733] = 18'b000000001111111100; 
assign wn_re[734] = 18'b000000000001011101; assign wn_im[734] = 18'b000000001111111011; 
assign wn_re[735] = 18'b000000000001100100; assign wn_im[735] = 18'b000000001111111011; 
assign wn_re[736] = 18'b000000000001101011; assign wn_im[736] = 18'b000000001111111010; 
assign wn_re[737] = 18'b000000000001110001; assign wn_im[737] = 18'b000000001111111001; 
assign wn_re[738] = 18'b000000000001111000; assign wn_im[738] = 18'b000000001111111000; 
assign wn_re[739] = 18'b000000000001111111; assign wn_im[739] = 18'b000000001111111000; 
assign wn_re[740] = 18'b000000000010000101; assign wn_im[740] = 18'b000000001111110111; 
assign wn_re[741] = 18'b000000000010001100; assign wn_im[741] = 18'b000000001111110110; 
assign wn_re[742] = 18'b000000000010010010; assign wn_im[742] = 18'b000000001111110101; 
assign wn_re[743] = 18'b000000000010011001; assign wn_im[743] = 18'b000000001111110100; 
assign wn_re[744] = 18'b000000000010100000; assign wn_im[744] = 18'b000000001111110011; 
assign wn_re[745] = 18'b000000000010100110; assign wn_im[745] = 18'b000000001111110010; 
assign wn_re[746] = 18'b000000000010101101; assign wn_im[746] = 18'b000000001111110001; 
assign wn_re[747] = 18'b000000000010110100; assign wn_im[747] = 18'b000000001111110000; 
assign wn_re[748] = 18'b000000000010111010; assign wn_im[748] = 18'b000000001111101110; 
assign wn_re[749] = 18'b000000000011000001; assign wn_im[749] = 18'b000000001111101101; 
assign wn_re[750] = 18'b000000000011000111; assign wn_im[750] = 18'b000000001111101100; 
assign wn_re[751] = 18'b000000000011001110; assign wn_im[751] = 18'b000000001111101010; 
assign wn_re[752] = 18'b000000000011010100; assign wn_im[752] = 18'b000000001111101001; 
assign wn_re[753] = 18'b000000000011011011; assign wn_im[753] = 18'b000000001111101000; 
assign wn_re[754] = 18'b000000000011100001; assign wn_im[754] = 18'b000000001111100110; 
assign wn_re[755] = 18'b000000000011101000; assign wn_im[755] = 18'b000000001111100101; 
assign wn_re[756] = 18'b000000000011101111; assign wn_im[756] = 18'b000000001111100011; 
assign wn_re[757] = 18'b000000000011110101; assign wn_im[757] = 18'b000000001111100010; 
assign wn_re[758] = 18'b000000000011111100; assign wn_im[758] = 18'b000000001111100000; 
assign wn_re[759] = 18'b000000000100000010; assign wn_im[759] = 18'b000000001111011110; 
assign wn_re[760] = 18'b000000000100001001; assign wn_im[760] = 18'b000000001111011101; 
assign wn_re[761] = 18'b000000000100001111; assign wn_im[761] = 18'b000000001111011011; 
assign wn_re[762] = 18'b000000000100010101; assign wn_im[762] = 18'b000000001111011001; 
assign wn_re[763] = 18'b000000000100011100; assign wn_im[763] = 18'b000000001111010111; 
assign wn_re[764] = 18'b000000000100100010; assign wn_im[764] = 18'b000000001111010101; 
assign wn_re[765] = 18'b000000000100101001; assign wn_im[765] = 18'b000000001111010011; 
assign wn_re[766] = 18'b000000000100101111; assign wn_im[766] = 18'b000000001111010001; 
assign wn_re[767] = 18'b000000000100110110; assign wn_im[767] = 18'b000000001111001111; 
assign wn_re[768] = 18'b000000000100111100; assign wn_im[768] = 18'b000000001111001101; 
assign wn_re[769] = 18'b000000000101000010; assign wn_im[769] = 18'b000000001111001011; 
assign wn_re[770] = 18'b000000000101001001; assign wn_im[770] = 18'b000000001111001001; 
assign wn_re[771] = 18'b000000000101001111; assign wn_im[771] = 18'b000000001111000111; 
assign wn_re[772] = 18'b000000000101010101; assign wn_im[772] = 18'b000000001111000101; 
assign wn_re[773] = 18'b000000000101011100; assign wn_im[773] = 18'b000000001111000011; 
assign wn_re[774] = 18'b000000000101100010; assign wn_im[774] = 18'b000000001111000000; 
assign wn_re[775] = 18'b000000000101101000; assign wn_im[775] = 18'b000000001110111110; 
assign wn_re[776] = 18'b000000000101101110; assign wn_im[776] = 18'b000000001110111011; 
assign wn_re[777] = 18'b000000000101110101; assign wn_im[777] = 18'b000000001110111001; 
assign wn_re[778] = 18'b000000000101111011; assign wn_im[778] = 18'b000000001110110111; 
assign wn_re[779] = 18'b000000000110000001; assign wn_im[779] = 18'b000000001110110100; 
assign wn_re[780] = 18'b000000000110000111; assign wn_im[780] = 18'b000000001110110010; 
assign wn_re[781] = 18'b000000000110001110; assign wn_im[781] = 18'b000000001110101111; 
assign wn_re[782] = 18'b000000000110010100; assign wn_im[782] = 18'b000000001110101100; 
assign wn_re[783] = 18'b000000000110011010; assign wn_im[783] = 18'b000000001110101010; 
assign wn_re[784] = 18'b000000000110100000; assign wn_im[784] = 18'b000000001110100111; 
assign wn_re[785] = 18'b000000000110100110; assign wn_im[785] = 18'b000000001110100100; 
assign wn_re[786] = 18'b000000000110101100; assign wn_im[786] = 18'b000000001110100001; 
assign wn_re[787] = 18'b000000000110110010; assign wn_im[787] = 18'b000000001110011111; 
assign wn_re[788] = 18'b000000000110111000; assign wn_im[788] = 18'b000000001110011100; 
assign wn_re[789] = 18'b000000000110111110; assign wn_im[789] = 18'b000000001110011001; 
assign wn_re[790] = 18'b000000000111000100; assign wn_im[790] = 18'b000000001110010110; 
assign wn_re[791] = 18'b000000000111001010; assign wn_im[791] = 18'b000000001110010011; 
assign wn_re[792] = 18'b000000000111010000; assign wn_im[792] = 18'b000000001110010000; 
assign wn_re[793] = 18'b000000000111010110; assign wn_im[793] = 18'b000000001110001101; 
assign wn_re[794] = 18'b000000000111011100; assign wn_im[794] = 18'b000000001110001010; 
assign wn_re[795] = 18'b000000000111100010; assign wn_im[795] = 18'b000000001110000111; 
assign wn_re[796] = 18'b000000000111101000; assign wn_im[796] = 18'b000000001110000011; 
assign wn_re[797] = 18'b000000000111101110; assign wn_im[797] = 18'b000000001110000000; 
assign wn_re[798] = 18'b000000000111110100; assign wn_im[798] = 18'b000000001101111101; 
assign wn_re[799] = 18'b000000000111111010; assign wn_im[799] = 18'b000000001101111010; 
assign wn_re[800] = 18'b000000001000000000; assign wn_im[800] = 18'b000000001101110110; 
assign wn_re[801] = 18'b000000001000000101; assign wn_im[801] = 18'b000000001101110011; 
assign wn_re[802] = 18'b000000001000001011; assign wn_im[802] = 18'b000000001101110000; 
assign wn_re[803] = 18'b000000001000010001; assign wn_im[803] = 18'b000000001101101100; 
assign wn_re[804] = 18'b000000001000010111; assign wn_im[804] = 18'b000000001101101001; 
assign wn_re[805] = 18'b000000001000011100; assign wn_im[805] = 18'b000000001101100101; 
assign wn_re[806] = 18'b000000001000100010; assign wn_im[806] = 18'b000000001101100010; 
assign wn_re[807] = 18'b000000001000101000; assign wn_im[807] = 18'b000000001101011110; 
assign wn_re[808] = 18'b000000001000101101; assign wn_im[808] = 18'b000000001101011010; 
assign wn_re[809] = 18'b000000001000110011; assign wn_im[809] = 18'b000000001101010111; 
assign wn_re[810] = 18'b000000001000111000; assign wn_im[810] = 18'b000000001101010011; 
assign wn_re[811] = 18'b000000001000111110; assign wn_im[811] = 18'b000000001101001111; 
assign wn_re[812] = 18'b000000001001000011; assign wn_im[812] = 18'b000000001101001011; 
assign wn_re[813] = 18'b000000001001001001; assign wn_im[813] = 18'b000000001101001000; 
assign wn_re[814] = 18'b000000001001001110; assign wn_im[814] = 18'b000000001101000100; 
assign wn_re[815] = 18'b000000001001010100; assign wn_im[815] = 18'b000000001101000000; 
assign wn_re[816] = 18'b000000001001011001; assign wn_im[816] = 18'b000000001100111100; 
assign wn_re[817] = 18'b000000001001011111; assign wn_im[817] = 18'b000000001100111000; 
assign wn_re[818] = 18'b000000001001100100; assign wn_im[818] = 18'b000000001100110100; 
assign wn_re[819] = 18'b000000001001101010; assign wn_im[819] = 18'b000000001100110000; 
assign wn_re[820] = 18'b000000001001101111; assign wn_im[820] = 18'b000000001100101100; 
assign wn_re[821] = 18'b000000001001110100; assign wn_im[821] = 18'b000000001100101000; 
assign wn_re[822] = 18'b000000001001111001; assign wn_im[822] = 18'b000000001100100100; 
assign wn_re[823] = 18'b000000001001111111; assign wn_im[823] = 18'b000000001100011111; 
assign wn_re[824] = 18'b000000001010000100; assign wn_im[824] = 18'b000000001100011011; 
assign wn_re[825] = 18'b000000001010001001; assign wn_im[825] = 18'b000000001100010111; 
assign wn_re[826] = 18'b000000001010001110; assign wn_im[826] = 18'b000000001100010011; 
assign wn_re[827] = 18'b000000001010010011; assign wn_im[827] = 18'b000000001100001110; 
assign wn_re[828] = 18'b000000001010011001; assign wn_im[828] = 18'b000000001100001010; 
assign wn_re[829] = 18'b000000001010011110; assign wn_im[829] = 18'b000000001100000110; 
assign wn_re[830] = 18'b000000001010100011; assign wn_im[830] = 18'b000000001100000001; 
assign wn_re[831] = 18'b000000001010101000; assign wn_im[831] = 18'b000000001011111101; 
assign wn_re[832] = 18'b000000001010101101; assign wn_im[832] = 18'b000000001011111000; 
assign wn_re[833] = 18'b000000001010110010; assign wn_im[833] = 18'b000000001011110100; 
assign wn_re[834] = 18'b000000001010110111; assign wn_im[834] = 18'b000000001011101111; 
assign wn_re[835] = 18'b000000001010111011; assign wn_im[835] = 18'b000000001011101011; 
assign wn_re[836] = 18'b000000001011000000; assign wn_im[836] = 18'b000000001011100110; 
assign wn_re[837] = 18'b000000001011000101; assign wn_im[837] = 18'b000000001011100010; 
assign wn_re[838] = 18'b000000001011001010; assign wn_im[838] = 18'b000000001011011101; 
assign wn_re[839] = 18'b000000001011001111; assign wn_im[839] = 18'b000000001011011000; 
assign wn_re[840] = 18'b000000001011010100; assign wn_im[840] = 18'b000000001011010100; 
assign wn_re[841] = 18'b000000001011011000; assign wn_im[841] = 18'b000000001011001111; 
assign wn_re[842] = 18'b000000001011011101; assign wn_im[842] = 18'b000000001011001010; 
assign wn_re[843] = 18'b000000001011100010; assign wn_im[843] = 18'b000000001011000101; 
assign wn_re[844] = 18'b000000001011100110; assign wn_im[844] = 18'b000000001011000000; 
assign wn_re[845] = 18'b000000001011101011; assign wn_im[845] = 18'b000000001010111011; 
assign wn_re[846] = 18'b000000001011101111; assign wn_im[846] = 18'b000000001010110111; 
assign wn_re[847] = 18'b000000001011110100; assign wn_im[847] = 18'b000000001010110010; 
assign wn_re[848] = 18'b000000001011111000; assign wn_im[848] = 18'b000000001010101101; 
assign wn_re[849] = 18'b000000001011111101; assign wn_im[849] = 18'b000000001010101000; 
assign wn_re[850] = 18'b000000001100000001; assign wn_im[850] = 18'b000000001010100011; 
assign wn_re[851] = 18'b000000001100000110; assign wn_im[851] = 18'b000000001010011110; 
assign wn_re[852] = 18'b000000001100001010; assign wn_im[852] = 18'b000000001010011001; 
assign wn_re[853] = 18'b000000001100001110; assign wn_im[853] = 18'b000000001010010011; 
assign wn_re[854] = 18'b000000001100010011; assign wn_im[854] = 18'b000000001010001110; 
assign wn_re[855] = 18'b000000001100010111; assign wn_im[855] = 18'b000000001010001001; 
assign wn_re[856] = 18'b000000001100011011; assign wn_im[856] = 18'b000000001010000100; 
assign wn_re[857] = 18'b000000001100011111; assign wn_im[857] = 18'b000000001001111111; 
assign wn_re[858] = 18'b000000001100100100; assign wn_im[858] = 18'b000000001001111001; 
assign wn_re[859] = 18'b000000001100101000; assign wn_im[859] = 18'b000000001001110100; 
assign wn_re[860] = 18'b000000001100101100; assign wn_im[860] = 18'b000000001001101111; 
assign wn_re[861] = 18'b000000001100110000; assign wn_im[861] = 18'b000000001001101010; 
assign wn_re[862] = 18'b000000001100110100; assign wn_im[862] = 18'b000000001001100100; 
assign wn_re[863] = 18'b000000001100111000; assign wn_im[863] = 18'b000000001001011111; 
assign wn_re[864] = 18'b000000001100111100; assign wn_im[864] = 18'b000000001001011001; 
assign wn_re[865] = 18'b000000001101000000; assign wn_im[865] = 18'b000000001001010100; 
assign wn_re[866] = 18'b000000001101000100; assign wn_im[866] = 18'b000000001001001110; 
assign wn_re[867] = 18'b000000001101001000; assign wn_im[867] = 18'b000000001001001001; 
assign wn_re[868] = 18'b000000001101001011; assign wn_im[868] = 18'b000000001001000011; 
assign wn_re[869] = 18'b000000001101001111; assign wn_im[869] = 18'b000000001000111110; 
assign wn_re[870] = 18'b000000001101010011; assign wn_im[870] = 18'b000000001000111000; 
assign wn_re[871] = 18'b000000001101010111; assign wn_im[871] = 18'b000000001000110011; 
assign wn_re[872] = 18'b000000001101011010; assign wn_im[872] = 18'b000000001000101101; 
assign wn_re[873] = 18'b000000001101011110; assign wn_im[873] = 18'b000000001000101000; 
assign wn_re[874] = 18'b000000001101100010; assign wn_im[874] = 18'b000000001000100010; 
assign wn_re[875] = 18'b000000001101100101; assign wn_im[875] = 18'b000000001000011100; 
assign wn_re[876] = 18'b000000001101101001; assign wn_im[876] = 18'b000000001000010111; 
assign wn_re[877] = 18'b000000001101101100; assign wn_im[877] = 18'b000000001000010001; 
assign wn_re[878] = 18'b000000001101110000; assign wn_im[878] = 18'b000000001000001011; 
assign wn_re[879] = 18'b000000001101110011; assign wn_im[879] = 18'b000000001000000101; 
assign wn_re[880] = 18'b000000001101110110; assign wn_im[880] = 18'b000000000111111111; 
assign wn_re[881] = 18'b000000001101111010; assign wn_im[881] = 18'b000000000111111010; 
assign wn_re[882] = 18'b000000001101111101; assign wn_im[882] = 18'b000000000111110100; 
assign wn_re[883] = 18'b000000001110000000; assign wn_im[883] = 18'b000000000111101110; 
assign wn_re[884] = 18'b000000001110000011; assign wn_im[884] = 18'b000000000111101000; 
assign wn_re[885] = 18'b000000001110000111; assign wn_im[885] = 18'b000000000111100010; 
assign wn_re[886] = 18'b000000001110001010; assign wn_im[886] = 18'b000000000111011100; 
assign wn_re[887] = 18'b000000001110001101; assign wn_im[887] = 18'b000000000111010110; 
assign wn_re[888] = 18'b000000001110010000; assign wn_im[888] = 18'b000000000111010000; 
assign wn_re[889] = 18'b000000001110010011; assign wn_im[889] = 18'b000000000111001010; 
assign wn_re[890] = 18'b000000001110010110; assign wn_im[890] = 18'b000000000111000100; 
assign wn_re[891] = 18'b000000001110011001; assign wn_im[891] = 18'b000000000110111110; 
assign wn_re[892] = 18'b000000001110011100; assign wn_im[892] = 18'b000000000110111000; 
assign wn_re[893] = 18'b000000001110011111; assign wn_im[893] = 18'b000000000110110010; 
assign wn_re[894] = 18'b000000001110100001; assign wn_im[894] = 18'b000000000110101100; 
assign wn_re[895] = 18'b000000001110100100; assign wn_im[895] = 18'b000000000110100110; 
assign wn_re[896] = 18'b000000001110100111; assign wn_im[896] = 18'b000000000110100000; 
assign wn_re[897] = 18'b000000001110101010; assign wn_im[897] = 18'b000000000110011010; 
assign wn_re[898] = 18'b000000001110101100; assign wn_im[898] = 18'b000000000110010100; 
assign wn_re[899] = 18'b000000001110101111; assign wn_im[899] = 18'b000000000110001110; 
assign wn_re[900] = 18'b000000001110110010; assign wn_im[900] = 18'b000000000110000111; 
assign wn_re[901] = 18'b000000001110110100; assign wn_im[901] = 18'b000000000110000001; 
assign wn_re[902] = 18'b000000001110110111; assign wn_im[902] = 18'b000000000101111011; 
assign wn_re[903] = 18'b000000001110111001; assign wn_im[903] = 18'b000000000101110101; 
assign wn_re[904] = 18'b000000001110111011; assign wn_im[904] = 18'b000000000101101110; 
assign wn_re[905] = 18'b000000001110111110; assign wn_im[905] = 18'b000000000101101000; 
assign wn_re[906] = 18'b000000001111000000; assign wn_im[906] = 18'b000000000101100010; 
assign wn_re[907] = 18'b000000001111000011; assign wn_im[907] = 18'b000000000101011100; 
assign wn_re[908] = 18'b000000001111000101; assign wn_im[908] = 18'b000000000101010101; 
assign wn_re[909] = 18'b000000001111000111; assign wn_im[909] = 18'b000000000101001111; 
assign wn_re[910] = 18'b000000001111001001; assign wn_im[910] = 18'b000000000101001001; 
assign wn_re[911] = 18'b000000001111001011; assign wn_im[911] = 18'b000000000101000010; 
assign wn_re[912] = 18'b000000001111001101; assign wn_im[912] = 18'b000000000100111100; 
assign wn_re[913] = 18'b000000001111001111; assign wn_im[913] = 18'b000000000100110110; 
assign wn_re[914] = 18'b000000001111010001; assign wn_im[914] = 18'b000000000100101111; 
assign wn_re[915] = 18'b000000001111010011; assign wn_im[915] = 18'b000000000100101001; 
assign wn_re[916] = 18'b000000001111010101; assign wn_im[916] = 18'b000000000100100010; 
assign wn_re[917] = 18'b000000001111010111; assign wn_im[917] = 18'b000000000100011100; 
assign wn_re[918] = 18'b000000001111011001; assign wn_im[918] = 18'b000000000100010101; 
assign wn_re[919] = 18'b000000001111011011; assign wn_im[919] = 18'b000000000100001111; 
assign wn_re[920] = 18'b000000001111011101; assign wn_im[920] = 18'b000000000100001001; 
assign wn_re[921] = 18'b000000001111011110; assign wn_im[921] = 18'b000000000100000010; 
assign wn_re[922] = 18'b000000001111100000; assign wn_im[922] = 18'b000000000011111100; 
assign wn_re[923] = 18'b000000001111100010; assign wn_im[923] = 18'b000000000011110101; 
assign wn_re[924] = 18'b000000001111100011; assign wn_im[924] = 18'b000000000011101111; 
assign wn_re[925] = 18'b000000001111100101; assign wn_im[925] = 18'b000000000011101000; 
assign wn_re[926] = 18'b000000001111100110; assign wn_im[926] = 18'b000000000011100001; 
assign wn_re[927] = 18'b000000001111101000; assign wn_im[927] = 18'b000000000011011011; 
assign wn_re[928] = 18'b000000001111101001; assign wn_im[928] = 18'b000000000011010100; 
assign wn_re[929] = 18'b000000001111101010; assign wn_im[929] = 18'b000000000011001110; 
assign wn_re[930] = 18'b000000001111101100; assign wn_im[930] = 18'b000000000011000111; 
assign wn_re[931] = 18'b000000001111101101; assign wn_im[931] = 18'b000000000011000001; 
assign wn_re[932] = 18'b000000001111101110; assign wn_im[932] = 18'b000000000010111010; 
assign wn_re[933] = 18'b000000001111110000; assign wn_im[933] = 18'b000000000010110100; 
assign wn_re[934] = 18'b000000001111110001; assign wn_im[934] = 18'b000000000010101101; 
assign wn_re[935] = 18'b000000001111110010; assign wn_im[935] = 18'b000000000010100110; 
assign wn_re[936] = 18'b000000001111110011; assign wn_im[936] = 18'b000000000010100000; 
assign wn_re[937] = 18'b000000001111110100; assign wn_im[937] = 18'b000000000010011001; 
assign wn_re[938] = 18'b000000001111110101; assign wn_im[938] = 18'b000000000010010010; 
assign wn_re[939] = 18'b000000001111110110; assign wn_im[939] = 18'b000000000010001100; 
assign wn_re[940] = 18'b000000001111110111; assign wn_im[940] = 18'b000000000010000101; 
assign wn_re[941] = 18'b000000001111111000; assign wn_im[941] = 18'b000000000001111111; 
assign wn_re[942] = 18'b000000001111111000; assign wn_im[942] = 18'b000000000001111000; 
assign wn_re[943] = 18'b000000001111111001; assign wn_im[943] = 18'b000000000001110001; 
assign wn_re[944] = 18'b000000001111111010; assign wn_im[944] = 18'b000000000001101011; 
assign wn_re[945] = 18'b000000001111111011; assign wn_im[945] = 18'b000000000001100100; 
assign wn_re[946] = 18'b000000001111111011; assign wn_im[946] = 18'b000000000001011101; 
assign wn_re[947] = 18'b000000001111111100; assign wn_im[947] = 18'b000000000001010111; 
assign wn_re[948] = 18'b000000001111111100; assign wn_im[948] = 18'b000000000001010000; 
assign wn_re[949] = 18'b000000001111111101; assign wn_im[949] = 18'b000000000001001001; 
assign wn_re[950] = 18'b000000001111111101; assign wn_im[950] = 18'b000000000001000010; 
assign wn_re[951] = 18'b000000001111111110; assign wn_im[951] = 18'b000000000000111100; 
assign wn_re[952] = 18'b000000001111111110; assign wn_im[952] = 18'b000000000000110101; 
assign wn_re[953] = 18'b000000001111111110; assign wn_im[953] = 18'b000000000000101110; 
assign wn_re[954] = 18'b000000001111111111; assign wn_im[954] = 18'b000000000000101000; 
assign wn_re[955] = 18'b000000001111111111; assign wn_im[955] = 18'b000000000000100001; 
assign wn_re[956] = 18'b000000001111111111; assign wn_im[956] = 18'b000000000000011010; 
assign wn_re[957] = 18'b000000001111111111; assign wn_im[957] = 18'b000000000000010100; 
assign wn_re[958] = 18'b000000001111111111; assign wn_im[958] = 18'b000000000000001101; 
assign wn_re[959] = 18'b000000001111111111; assign wn_im[959] = 18'b000000000000000110; 

endmodule
